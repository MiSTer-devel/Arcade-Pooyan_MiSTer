library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity pooyan_char_grphx1 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(11 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of pooyan_char_grphx1 is
	type rom is array(0 to  4095) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"30",X"30",X"30",X"10",X"10",X"00",X"00",X"00",X"00",X"00",X"80",X"C0",X"F0",X"F0",X"30",X"00",
		X"00",X"10",X"30",X"00",X"F0",X"F0",X"F0",X"00",X"C0",X"80",X"00",X"00",X"C0",X"E0",X"C0",X"00",
		X"00",X"00",X"00",X"00",X"30",X"30",X"10",X"00",X"00",X"10",X"10",X"70",X"F0",X"E0",X"C0",X"00",
		X"F0",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"00",X"33",X"33",X"CC",X"19",
		X"00",X"88",X"44",X"00",X"00",X"55",X"22",X"00",X"30",X"33",X"30",X"30",X"33",X"30",X"20",X"00",
		X"13",X"13",X"13",X"03",X"00",X"00",X"00",X"00",X"0F",X"0F",X"09",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"F0",X"F0",X"FF",X"F0",X"F0",X"FF",X"F0",X"CC",X"C0",X"C0",X"CC",X"C0",X"C0",X"CC",X"C0",
		X"FF",X"EE",X"BB",X"22",X"22",X"55",X"30",X"70",X"88",X"11",X"00",X"40",X"C0",X"CC",X"C0",X"C0",
		X"F0",X"FF",X"E0",X"C0",X"88",X"44",X"EE",X"00",X"80",X"44",X"44",X"00",X"00",X"00",X"00",X"00",
		X"00",X"88",X"F9",X"FF",X"F9",X"F9",X"F9",X"88",X"30",X"33",X"E2",X"E2",X"E2",X"EE",X"E2",X"00",
		X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0C",X"0C",X"0C",X"0C",X"0F",X"0F",X"0F",X"00",X"00",X"02",X"06",X"0C",X"0C",X"08",X"00",X"00",
		X"0C",X"0C",X"04",X"0C",X"0C",X"04",X"0C",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"51",X"31",X"50",X"75",X"00",X"00",X"33",X"FF",X"FF",X"FF",X"FF",X"FE",
		X"00",X"10",X"60",X"30",X"00",X"00",X"00",X"00",X"F0",X"F7",X"77",X"F0",X"F1",X"00",X"00",X"00",
		X"00",X"01",X"01",X"70",X"F0",X"D0",X"00",X"00",X"0C",X"08",X"68",X"24",X"E0",X"60",X"08",X"0C",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"CC",X"00",X"00",X"88",X"88",X"88",X"88",X"00",X"00",X"00",X"11",X"23",X"11",X"00",X"00",X"00",
		X"77",X"77",X"77",X"33",X"51",X"00",X"00",X"00",X"FE",X"FE",X"FF",X"FF",X"FF",X"FF",X"33",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"55",X"11",X"00",X"22",X"00",X"00",X"00",X"88",X"EE",X"FF",
		X"00",X"0F",X"01",X"CC",X"FF",X"00",X"11",X"CC",X"17",X"3F",X"3F",X"37",X"FF",X"00",X"EE",X"FF",
		X"00",X"00",X"00",X"70",X"F0",X"D0",X"00",X"00",X"06",X"0E",X"2C",X"24",X"E0",X"60",X"0C",X"06",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"33",X"76",X"33",X"03",X"01",X"13",X"BB",X"EE",X"99",X"DD",X"9B",X"07",X"CF",X"DF",X"FF",X"11",
		X"00",X"77",X"11",X"00",X"00",X"08",X"08",X"04",X"00",X"00",X"88",X"44",X"22",X"00",X"00",X"04",
		X"11",X"22",X"CC",X"33",X"00",X"0C",X"0F",X"07",X"88",X"44",X"00",X"00",X"00",X"07",X"0F",X"08",
		X"00",X"11",X"66",X"88",X"00",X"13",X"67",X"88",X"66",X"99",X"00",X"00",X"00",X"08",X"00",X"00",
		X"33",X"22",X"CC",X"00",X"00",X"11",X"EE",X"00",X"88",X"00",X"00",X"33",X"44",X"88",X"00",X"00",
		X"00",X"00",X"00",X"FF",X"FF",X"88",X"00",X"00",X"00",X"00",X"FF",X"FF",X"88",X"00",X"00",X"00",
		X"00",X"AA",X"22",X"11",X"00",X"00",X"88",X"00",X"00",X"00",X"CC",X"66",X"11",X"EE",X"66",X"11",
		X"66",X"26",X"33",X"00",X"00",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"33",X"CC",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"CC",X"22",X"11",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"CC",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"33",X"88",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"1F",X"BF",X"FE",X"A8",X"60",X"C0",X"80",X"00",X"C0",X"C0",X"51",X"31",X"11",X"00",X"00",X"00",
		X"00",X"11",X"33",X"47",X"8C",X"01",X"33",X"00",X"33",X"FF",X"CC",X"00",X"00",X"0E",X"FF",X"33",
		X"33",X"46",X"8C",X"00",X"00",X"11",X"33",X"33",X"00",X"00",X"00",X"00",X"33",X"FF",X"EE",X"88",
		X"3F",X"37",X"3F",X"13",X"13",X"3F",X"37",X"3F",X"8C",X"CE",X"CF",X"8F",X"8E",X"CE",X"CC",X"8C",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0C",X"26",X"17",X"13",X"13",X"13",X"01",X"00",X"00",X"00",X"88",X"88",X"CC",X"CC",X"EE",X"EE",
		X"CC",X"CC",X"6E",X"3F",X"DF",X"7F",X"7F",X"0F",X"00",X"00",X"00",X"88",X"88",X"CC",X"EE",X"6E",
		X"66",X"66",X"33",X"11",X"00",X"11",X"33",X"67",X"11",X"22",X"99",X"EE",X"3B",X"2A",X"7F",X"99",
		X"00",X"00",X"00",X"11",X"B3",X"73",X"B1",X"73",X"00",X"00",X"77",X"FF",X"FF",X"FF",X"FE",X"EC",
		X"00",X"11",X"33",X"37",X"13",X"13",X"00",X"00",X"88",X"88",X"00",X"00",X"88",X"0C",X"8C",X"00",
		X"00",X"00",X"00",X"23",X"23",X"11",X"00",X"00",X"00",X"00",X"02",X"00",X"08",X"0C",X"00",X"00",
		X"00",X"00",X"00",X"00",X"11",X"03",X"66",X"CC",X"00",X"00",X"00",X"00",X"08",X"00",X"00",X"00",
		X"33",X"33",X"01",X"01",X"01",X"00",X"00",X"00",X"6E",X"6E",X"6E",X"FF",X"6E",X"2E",X"2E",X"3F",
		X"DF",X"57",X"57",X"57",X"47",X"47",X"23",X"33",X"CC",X"CC",X"CC",X"EE",X"CC",X"CC",X"4C",X"4C",
		X"00",X"13",X"22",X"22",X"02",X"01",X"01",X"00",X"66",X"66",X"CC",X"CC",X"CC",X"66",X"66",X"66",
		X"CC",X"00",X"00",X"22",X"CC",X"11",X"00",X"11",X"04",X"00",X"DD",X"DD",X"BB",X"33",X"66",X"CC",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"BF",X"9F",X"07",X"03",X"06",X"08",X"00",X"13",X"9F",X"CE",X"CC",X"6E",X"66",X"33",X"00",
		X"04",X"04",X"08",X"09",X"09",X"1D",X"03",X"00",X"17",X"1F",X"3F",X"7F",X"EE",X"89",X"02",X"0C",
		X"00",X"00",X"00",X"00",X"88",X"CC",X"EF",X"3F",X"37",X"17",X"88",X"88",X"00",X"00",X"33",X"CF",
		X"00",X"00",X"00",X"88",X"CC",X"77",X"33",X"00",X"00",X"00",X"00",X"00",X"00",X"44",X"FF",X"BB",
		X"CC",X"89",X"13",X"1B",X"26",X"00",X"9B",X"45",X"19",X"2A",X"AA",X"AB",X"AB",X"CE",X"8C",X"08",
		X"EF",X"EF",X"4D",X"11",X"33",X"66",X"88",X"CC",X"89",X"CD",X"CD",X"BB",X"BB",X"33",X"11",X"11",
		X"44",X"44",X"44",X"44",X"88",X"00",X"00",X"88",X"00",X"00",X"00",X"00",X"00",X"CC",X"EE",X"33",
		X"44",X"23",X"0B",X"00",X"04",X"01",X"01",X"03",X"00",X"0F",X"00",X"00",X"00",X"0F",X"00",X"00",
		X"70",X"30",X"11",X"00",X"00",X"00",X"00",X"00",X"C0",X"C0",X"CC",X"C0",X"40",X"00",X"00",X"00",
		X"8B",X"01",X"44",X"47",X"03",X"03",X"02",X"01",X"00",X"0F",X"00",X"00",X"00",X"0F",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0E",X"07",X"8B",X"03",X"11",X"01",X"02",X"01",X"00",X"0F",X"00",X"00",X"00",X"0F",X"88",X"CC",
		X"00",X"00",X"20",X"50",X"20",X"50",X"20",X"00",X"00",X"44",X"33",X"11",X"FF",X"33",X"66",X"44",
		X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"33",X"CC",
		X"00",X"99",X"66",X"00",X"00",X"00",X"00",X"00",X"EE",X"00",X"EE",X"22",X"11",X"00",X"00",X"00",
		X"21",X"31",X"D1",X"70",X"10",X"00",X"22",X"76",X"0F",X"8F",X"F7",X"F2",X"F0",X"00",X"10",X"F0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"0F",X"0F",X"0F",X"0F",X"03",X"03",X"00",X"00",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"0F",X"1F",X"0F",X"1F",X"FF",X"4F",X"EF",X"8F",X"BF",X"EF",X"8F",X"CF",X"8F",X"8F",X"0F",X"0F",
		X"FF",X"FF",X"FF",X"EF",X"CF",X"FF",X"AF",X"1F",X"6F",X"5F",X"9F",X"FF",X"BF",X"FF",X"BF",X"7F",
		X"0F",X"6F",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",X"0F",X"0F",X"0F",X"4F",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"BF",X"0F",X"0F",X"0F",X"0F",X"EF",X"CF",X"8F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"00",X"00",X"00",X"00",X"00",X"06",X"0F",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"1F",X"1F",X"0F",X"0F",X"0F",X"1F",X"3F",X"BF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"01",X"FF",X"33",X"77",X"22",X"08",X"0D",X"0F",X"0F",
		X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"0F",X"0F",X"07",X"07",X"0F",X"0F",X"07",
		X"00",X"00",X"88",X"CC",X"CC",X"EE",X"E2",X"22",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"1F",X"2F",X"3F",X"1F",X"1F",X"3F",X"6F",X"3F",
		X"00",X"00",X"00",X"01",X"07",X"8F",X"CF",X"CF",X"00",X"60",X"F0",X"3C",X"0F",X"0F",X"0F",X"0F",
		X"00",X"B0",X"F0",X"F0",X"E1",X"0F",X"0F",X"0F",X"CF",X"78",X"E1",X"6D",X"ED",X"EF",X"6F",X"0F",
		X"0F",X"0F",X"07",X"03",X"07",X"0F",X"0F",X"07",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"00",X"00",X"00",X"00",X"80",X"E0",X"F0",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"C0",
		X"EE",X"7F",X"5F",X"9F",X"3F",X"6F",X"0F",X"1F",X"00",X"00",X"CC",X"CC",X"88",X"CC",X"EE",X"EE",
		X"88",X"CC",X"4C",X"88",X"EE",X"FF",X"7F",X"6E",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"F0",X"F0",X"C0",X"00",X"00",X"01",X"00",X"00",X"C0",X"F0",X"70",X"16",X"0F",X"7E",
		X"00",X"10",X"10",X"70",X"F0",X"C3",X"C3",X"87",X"C3",X"C3",X"87",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"10",X"30",X"30",X"21",X"61",X"43",X"43",
		X"88",X"CC",X"CC",X"EE",X"BF",X"0F",X"0F",X"0F",X"00",X"00",X"00",X"00",X"00",X"66",X"AE",X"1F",
		X"2F",X"6F",X"FF",X"7F",X"6E",X"FF",X"2F",X"0F",X"7F",X"EE",X"DD",X"44",X"00",X"88",X"EE",X"DF",
		X"0F",X"1F",X"0F",X"2F",X"3F",X"FF",X"FF",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"3F",X"FF",X"FF",X"FF",X"FF",X"BF",X"0F",X"0F",X"BF",X"FF",X"FF",X"FF",X"7F",X"2F",X"0F",X"0F",
		X"3F",X"7F",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",X"3F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"6E",X"BF",X"1F",X"3F",X"DD",X"88",X"33",X"FF",X"00",X"00",X"88",X"88",X"88",X"77",X"FF",X"FF",
		X"00",X"00",X"80",X"F0",X"F0",X"1E",X"0F",X"0F",X"00",X"00",X"F0",X"F0",X"F0",X"87",X"0F",X"0F",
		X"FF",X"FF",X"7F",X"FF",X"1F",X"7F",X"1F",X"3F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"0F",X"0F",X"0F",X"0F",X"06",X"00",X"00",X"00",X"0F",X"0F",X"0F",X"08",X"00",X"00",X"00",X"00",
		X"00",X"CC",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"88",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"F0",X"F0",X"E1",X"0F",X"0F",X"0F",X"0F",X"F0",X"F0",X"F0",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"0F",X"0F",X"08",X"00",X"00",X"00",X"00",X"00",X"0F",X"0F",X"03",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"CC",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"33",X"FF",X"FF",X"FF",X"FF",
		X"0F",X"0F",X"0F",X"0F",X"07",X"03",X"00",X"01",X"0F",X"0F",X"EF",X"6F",X"7F",X"7F",X"6E",X"CC",
		X"00",X"01",X"C1",X"F0",X"E1",X"0F",X"0E",X"19",X"0E",X"0F",X"0F",X"3F",X"1F",X"3F",X"6F",X"CF",
		X"0F",X"1F",X"2F",X"0F",X"0F",X"1F",X"0F",X"0F",X"6E",X"FF",X"7F",X"FF",X"EE",X"FF",X"7F",X"EE",
		X"8F",X"CF",X"67",X"33",X"67",X"67",X"CF",X"07",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"FF",X"7F",X"9F",X"3F",X"1F",X"7F",X"3F",X"0F",
		X"F0",X"F0",X"3C",X"0F",X"0F",X"0F",X"0F",X"0F",X"F0",X"E1",X"E1",X"C3",X"0F",X"0F",X"0F",X"0F",
		X"CF",X"EF",X"EE",X"FF",X"FF",X"FF",X"FF",X"FF",X"0F",X"0F",X"07",X"00",X"00",X"00",X"88",X"FF",
		X"00",X"00",X"C0",X"C0",X"80",X"80",X"00",X"00",X"20",X"20",X"00",X"00",X"40",X"80",X"00",X"00",
		X"52",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1E",X"1E",X"02",X"01",X"00",X"20",X"01",X"00",
		X"1E",X"2C",X"48",X"48",X"0C",X"08",X"00",X"00",X"86",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"0A",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"0A",X"0F",
		X"00",X"30",X"70",X"70",X"30",X"10",X"00",X"00",X"70",X"C0",X"00",X"80",X"F0",X"F0",X"70",X"00",
		X"00",X"00",X"00",X"10",X"F0",X"F0",X"E0",X"00",X"00",X"20",X"60",X"E0",X"C0",X"80",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"30",X"00",X"00",X"22",X"10",X"10",X"20",X"F0",X"F0",
		X"00",X"00",X"30",X"20",X"A0",X"B0",X"F0",X"F0",X"88",X"88",X"AA",X"22",X"44",X"88",X"11",X"71",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"20",X"40",X"73",X"40",X"20",X"10",
		X"10",X"C0",X"A8",X"98",X"F6",X"98",X"A8",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"10",X"20",X"31",X"20",X"10",X"00",X"60",X"E0",X"54",X"44",X"FB",X"44",X"54",
		X"00",X"00",X"00",X"00",X"80",X"80",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"20",X"51",X"40",X"51",X"20",X"10",
		X"10",X"D0",X"20",X"54",X"90",X"54",X"20",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"10",X"20",X"20",X"20",X"10",X"10",X"20",X"E0",X"10",X"AA",X"40",X"AA",X"10",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"B3",X"F7",X"76",X"76",X"76",X"F7",X"B3",X"00",X"88",X"C4",X"40",X"C0",X"40",X"C4",X"88",
		X"00",X"22",X"11",X"00",X"00",X"00",X"11",X"22",X"00",X"00",X"40",X"98",X"11",X"98",X"40",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"E0",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"C0",X"00",X"00",X"F0",X"F0",X"F0",X"F0",X"F0",X"30",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"E0",X"F0",X"F0",X"F0",X"F0",X"F0",X"E0",
		X"00",X"00",X"80",X"E0",X"F0",X"C0",X"00",X"00",X"00",X"00",X"10",X"70",X"F0",X"30",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"C0",X"C0",X"C0",X"C0",X"C0",X"E0",X"E0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"00",X"00",
		X"00",X"C0",X"F0",X"F0",X"F0",X"F0",X"00",X"00",X"00",X"30",X"F0",X"F0",X"F0",X"F0",X"00",X"00",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"0F",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"0F",X"00",X"00",
		X"FF",X"FF",X"FF",X"77",X"B3",X"11",X"00",X"00",X"FC",X"EC",X"FE",X"FF",X"FF",X"FF",X"77",X"00",
		X"0F",X"0A",X"0F",X"0A",X"0A",X"0F",X"0A",X"0F",X"0F",X"0A",X"0F",X"0A",X"0A",X"0F",X"0A",X"0F",
		X"E2",X"22",X"E2",X"EE",X"CC",X"CC",X"88",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"E4",X"64",X"E4",X"CC",X"88",X"88",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"88",X"88",X"CC",X"E4",X"64",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"80",X"C0",X"F0",X"F0",X"F0",X"F0",X"E0",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"01",X"00",X"00",X"00",X"00",X"0F",X"0F",X"0C",X"78",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"07",X"07",X"07",X"01",
		X"00",X"00",X"08",X"08",X"0C",X"0C",X"0F",X"0F",X"30",X"10",X"10",X"00",X"00",X"00",X"00",X"0E",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"30",X"30",X"00",X"00",X"00",X"00",X"00",
		X"E1",X"F0",X"F0",X"F0",X"30",X"00",X"00",X"00",X"1E",X"F0",X"F0",X"96",X"C3",X"F0",X"30",X"00",
		X"88",X"88",X"88",X"22",X"00",X"11",X"00",X"00",X"AA",X"54",X"30",X"33",X"30",X"30",X"33",X"30",
		X"F0",X"F0",X"F0",X"F0",X"30",X"00",X"00",X"00",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"60",X"00",
		X"C0",X"F0",X"F2",X"FC",X"EC",X"98",X"00",X"00",X"C4",X"C0",X"D1",X"31",X"11",X"C4",X"44",X"00",
		X"00",X"00",X"00",X"00",X"01",X"01",X"01",X"00",X"00",X"00",X"00",X"0F",X"0F",X"0C",X"78",X"34",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"07",X"0F",X"0F",X"07",X"07",X"70",X"F0",
		X"00",X"00",X"08",X"08",X"0C",X"0C",X"86",X"E1",X"30",X"30",X"30",X"10",X"00",X"00",X"00",X"68",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"30",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F0",X"F0",X"C3",X"21",X"10",X"00",X"00",X"00",X"F0",X"F0",X"F0",X"C3",X"5A",X"F0",X"30",X"00",
		X"00",X"00",X"0B",X"40",X"80",X"20",X"F0",X"F0",X"00",X"00",X"08",X"0C",X"06",X"02",X"02",X"83",
		X"F0",X"F0",X"F0",X"70",X"10",X"00",X"00",X"00",X"81",X"E1",X"F0",X"F0",X"F0",X"F0",X"60",X"20",
		X"00",X"0F",X"00",X"00",X"51",X"0F",X"50",X"75",X"00",X"0F",X"33",X"FF",X"FF",X"0F",X"FF",X"FE",
		X"00",X"0F",X"88",X"CC",X"CC",X"0F",X"F2",X"32",X"00",X"0F",X"00",X"60",X"F1",X"0F",X"F1",X"E0",
		X"77",X"0F",X"77",X"33",X"51",X"0F",X"00",X"00",X"FE",X"0F",X"FF",X"FF",X"FF",X"0F",X"33",X"00",
		X"F2",X"0F",X"F2",X"EE",X"CC",X"0F",X"88",X"00",X"E0",X"0F",X"F1",X"F1",X"F1",X"0F",X"00",X"00",
		X"00",X"0F",X"00",X"11",X"B3",X"0F",X"B1",X"FB",X"00",X"0F",X"77",X"FF",X"FF",X"0F",X"FC",X"C8",
		X"00",X"0F",X"00",X"88",X"98",X"0F",X"FC",X"FC",X"00",X"0F",X"22",X"E2",X"E2",X"0F",X"C0",X"C0",
		X"FF",X"0F",X"FF",X"77",X"B3",X"0F",X"00",X"00",X"F8",X"0F",X"FC",X"FF",X"FF",X"0F",X"77",X"00",
		X"FC",X"0F",X"FC",X"DC",X"98",X"0F",X"00",X"00",X"C0",X"0F",X"C0",X"C0",X"E2",X"0F",X"22",X"00",
		X"00",X"31",X"20",X"71",X"E0",X"71",X"70",X"30",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"00",
		X"00",X"00",X"CC",X"66",X"EE",X"44",X"EE",X"DC",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"10",X"31",X"31",X"F0",X"73",X"30",X"00",X"00",X"F3",X"FF",X"FE",X"F0",X"F0",X"F0",X"F0",X"30",
		X"EE",X"FE",X"FC",X"F1",X"F0",X"F0",X"80",X"00",X"80",X"91",X"DD",X"F9",X"D1",X"80",X"00",X"00",
		X"00",X"00",X"31",X"20",X"31",X"70",X"70",X"70",X"00",X"00",X"44",X"FF",X"77",X"66",X"AA",X"77",
		X"CC",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"30",X"30",X"71",X"31",X"70",X"F0",X"00",X"00",X"B3",X"F3",X"FF",X"FE",X"F0",X"F0",X"B0",X"00",
		X"73",X"FB",X"F8",X"F8",X"F0",X"80",X"00",X"00",X"88",X"CC",X"CC",X"D1",X"B1",X"C0",X"71",X"77",
		X"C0",X"60",X"FC",X"F2",X"F0",X"F0",X"F0",X"F0",X"00",X"11",X"71",X"51",X"C0",X"C0",X"C0",X"F3",
		X"00",X"00",X"30",X"A8",X"A0",X"F0",X"F0",X"F0",X"00",X"88",X"88",X"11",X"31",X"D1",X"80",X"80",
		X"F0",X"F0",X"F0",X"E0",X"E2",X"CC",X"00",X"00",X"E0",X"E0",X"F0",X"80",X"80",X"E2",X"22",X"00",
		X"F0",X"F0",X"F0",X"F0",X"D8",X"D0",X"80",X"00",X"EE",X"33",X"11",X"22",X"44",X"C4",X"44",X"00",
		X"00",X"00",X"00",X"11",X"F3",X"73",X"FF",X"FF",X"00",X"00",X"00",X"EE",X"FF",X"FF",X"FF",X"FF",
		X"10",X"10",X"00",X"00",X"00",X"88",X"88",X"8A",X"00",X"00",X"00",X"00",X"23",X"23",X"00",X"23",
		X"FF",X"FF",X"77",X"77",X"33",X"11",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FE",X"FF",X"E0",X"00",
		X"8B",X"89",X"CD",X"CC",X"98",X"10",X"00",X"00",X"23",X"01",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"91",X"F3",X"73",X"FF",X"FF",X"FF",X"00",X"00",X"EE",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"10",X"10",X"00",X"00",X"00",X"88",X"8A",X"8F",X"00",X"00",X"00",X"00",X"00",X"23",X"23",X"00",
		X"FF",X"77",X"77",X"33",X"11",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"70",X"00",X"00",
		X"89",X"CC",X"C4",X"89",X"10",X"10",X"00",X"00",X"23",X"23",X"01",X"00",X"00",X"00",X"00",X"00",
		X"11",X"F3",X"73",X"FF",X"FF",X"FF",X"FF",X"77",X"EE",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"10",X"10",X"88",X"88",X"8A",X"CF",X"CD",X"CC",X"00",X"00",X"00",X"00",X"00",X"22",X"23",X"01",
		X"77",X"33",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"70",X"00",X"00",X"00",X"00",
		X"C8",X"80",X"88",X"01",X"10",X"10",X"00",X"00",X"44",X"67",X"23",X"01",X"00",X"00",X"00",X"00",
		X"1E",X"2C",X"48",X"48",X"0C",X"08",X"00",X"00",X"86",X"D1",X"33",X"11",X"30",X"70",X"70",X"70",
		X"52",X"88",X"CC",X"88",X"C0",X"E0",X"E0",X"E0",X"1E",X"1E",X"02",X"01",X"00",X"20",X"01",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"30",X"70",X"70",X"70",X"30",X"11",X"33",X"11",
		X"C0",X"E0",X"E0",X"E0",X"C0",X"88",X"CC",X"88",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"30",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"70",X"F0",X"30",X"10",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"30",X"10",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"30",X"F0",X"70",X"10",X"00",X"11",X"33",
		X"00",X"00",X"00",X"00",X"10",X"30",X"00",X"00",X"FC",X"44",X"00",X"70",X"F0",X"F0",X"F0",X"70",
		X"00",X"00",X"00",X"10",X"70",X"F0",X"30",X"10",X"00",X"00",X"33",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"00",X"00",X"30",X"10",X"00",X"00",X"00",X"00",X"70",X"F0",X"F0",X"F0",X"70",X"00",X"00",X"00",
		X"10",X"30",X"F0",X"70",X"10",X"00",X"11",X"33",X"F0",X"F0",X"F0",X"F0",X"F0",X"33",X"10",X"F0",
		X"74",X"CC",X"00",X"70",X"F0",X"F0",X"F0",X"70",X"C0",X"60",X"FC",X"F2",X"F0",X"F0",X"F0",X"F0",
		X"00",X"00",X"33",X"F0",X"F0",X"F0",X"F0",X"F0",X"00",X"00",X"30",X"A8",X"E0",X"F0",X"F0",X"F0",
		X"70",X"F0",X"F0",X"F0",X"70",X"00",X"00",X"00",X"F0",X"F0",X"F0",X"E0",X"E2",X"CC",X"00",X"00",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"33",X"30",X"E0",X"F0",X"F0",X"F0",X"F0",X"D8",X"D0",X"80",X"00");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
