library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity pooyan_prog is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(14 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of pooyan_prog is
	type rom is array(0 to  32767) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"AF",X"32",X"80",X"A1",X"C3",X"92",X"00",X"FF",X"77",X"3C",X"23",X"77",X"3C",X"19",X"C9",X"FF",
		X"77",X"23",X"10",X"FC",X"C9",X"FF",X"FF",X"FF",X"77",X"23",X"10",X"FC",X"0D",X"20",X"F9",X"C9",
		X"85",X"6F",X"3E",X"00",X"8C",X"67",X"7E",X"C9",X"87",X"E1",X"5F",X"16",X"00",X"19",X"5E",X"23",
		X"56",X"EB",X"E9",X"FF",X"FF",X"FF",X"FF",X"FF",X"E5",X"26",X"88",X"3A",X"A0",X"88",X"6F",X"CB",
		X"7E",X"28",X"0E",X"72",X"2C",X"73",X"2C",X"7D",X"FE",X"C0",X"30",X"02",X"3E",X"C0",X"32",X"A0",
		X"88",X"E1",X"C9",X"0F",X"33",X"31",X"24",X"22",X"21",X"15",X"13",X"11",X"07",X"06",X"05",X"04",
		X"03",X"02",X"01",X"FF",X"FF",X"FF",X"C3",X"6D",X"06",X"00",X"11",X"22",X"04",X"31",X"06",X"15",
		X"02",X"33",X"07",X"21",X"03",X"24",X"05",X"13",X"01",X"00",X"33",X"05",X"61",X"BE",X"05",X"66",
		X"07",X"06",X"DD",X"A8",X"05",X"60",X"BC",X"04",X"A6",X"51",X"05",X"38",X"8A",X"06",X"AD",X"BA",
		X"05",X"CA",X"32",X"00",X"A0",X"31",X"00",X"90",X"32",X"00",X"88",X"06",X"08",X"C5",X"21",X"00",
		X"00",X"DD",X"21",X"79",X"00",X"11",X"00",X"00",X"4A",X"7B",X"86",X"5F",X"30",X"04",X"14",X"20",
		X"01",X"0C",X"2C",X"20",X"F4",X"24",X"7C",X"E6",X"0F",X"20",X"EE",X"32",X"00",X"A0",X"7B",X"DD",
		X"BE",X"00",X"20",X"0C",X"7A",X"DD",X"BE",X"01",X"20",X"06",X"79",X"DD",X"BE",X"02",X"28",X"02",
		X"18",X"06",X"E5",X"21",X"FF",X"8F",X"34",X"E1",X"DD",X"23",X"DD",X"23",X"DD",X"23",X"10",X"C5",
		X"3A",X"E0",X"A0",X"E6",X"0F",X"21",X"69",X"00",X"E7",X"7E",X"B7",X"18",X"16",X"57",X"E6",X"0F",
		X"5F",X"AA",X"0F",X"0F",X"0F",X"0F",X"CD",X"FA",X"00",X"7B",X"FE",X"0A",X"38",X"02",X"C6",X"07",
		X"77",X"09",X"C9",X"32",X"00",X"A0",X"21",X"00",X"88",X"11",X"01",X"88",X"01",X"FD",X"07",X"36",
		X"00",X"ED",X"B0",X"3E",X"08",X"32",X"42",X"8A",X"21",X"C0",X"88",X"06",X"40",X"3E",X"FF",X"D7",
		X"21",X"43",X"8A",X"06",X"1C",X"D7",X"21",X"43",X"43",X"22",X"40",X"8A",X"32",X"00",X"A0",X"3E",
		X"01",X"32",X"87",X"A1",X"32",X"1F",X"88",X"21",X"C0",X"C0",X"22",X"A0",X"88",X"21",X"00",X"80",
		X"11",X"01",X"80",X"36",X"10",X"01",X"00",X"04",X"ED",X"B0",X"CD",X"E6",X"02",X"32",X"00",X"A0",
		X"3A",X"00",X"A0",X"2F",X"0F",X"0F",X"47",X"E6",X"01",X"32",X"0F",X"88",X"78",X"0F",X"47",X"E6",
		X"01",X"32",X"00",X"88",X"78",X"0F",X"47",X"E6",X"07",X"32",X"20",X"88",X"78",X"0F",X"0F",X"0F",
		X"47",X"E6",X"01",X"32",X"21",X"88",X"3A",X"00",X"A0",X"2F",X"E6",X"03",X"FE",X"03",X"28",X"04",
		X"C6",X"03",X"18",X"02",X"3E",X"FF",X"32",X"07",X"88",X"3A",X"E0",X"A0",X"47",X"E6",X"F0",X"0F",
		X"0F",X"0F",X"0F",X"21",X"53",X"00",X"E7",X"32",X"2F",X"88",X"78",X"E6",X"0F",X"21",X"53",X"00",
		X"E7",X"32",X"2C",X"88",X"32",X"00",X"A0",X"CD",X"EA",X"01",X"AF",X"CD",X"8F",X"0E",X"3E",X"01",
		X"32",X"80",X"A1",X"21",X"00",X"8A",X"06",X"0A",X"36",X"00",X"2C",X"36",X"00",X"2C",X"36",X"01",
		X"2C",X"10",X"F5",X"21",X"AA",X"88",X"36",X"01",X"32",X"00",X"A0",X"21",X"C0",X"89",X"AF",X"06",
		X"1E",X"D7",X"C3",X"0F",X"02",X"32",X"00",X"A0",X"18",X"FB",X"0B",X"32",X"00",X"A0",X"3A",X"80",
		X"A0",X"CB",X"5F",X"C0",X"78",X"B1",X"20",X"F2",X"37",X"C9",X"21",X"10",X"94",X"06",X"30",X"D7",
		X"21",X"10",X"90",X"06",X"30",X"D7",X"21",X"40",X"84",X"11",X"41",X"84",X"01",X"BF",X"03",X"36",
		X"1E",X"ED",X"B0",X"00",X"00",X"00",X"10",X"FB",X"32",X"00",X"A0",X"0D",X"20",X"F5",X"C9",X"26",
		X"88",X"3A",X"A1",X"88",X"6F",X"7E",X"87",X"30",X"05",X"CD",X"54",X"02",X"18",X"F1",X"E6",X"1F",
		X"4F",X"06",X"00",X"36",X"FF",X"23",X"5E",X"36",X"FF",X"2C",X"7D",X"FE",X"C0",X"30",X"02",X"3E",
		X"C0",X"32",X"A1",X"88",X"7B",X"21",X"42",X"02",X"09",X"5E",X"23",X"56",X"21",X"0F",X"02",X"E5",
		X"EB",X"E9",X"9B",X"03",X"C2",X"03",X"E9",X"03",X"96",X"04",X"52",X"05",X"6B",X"05",X"B2",X"05",
		X"EE",X"05",X"44",X"06",X"3A",X"3F",X"88",X"47",X"E6",X"0F",X"CA",X"61",X"02",X"CD",X"8C",X"20",
		X"C9",X"3A",X"06",X"88",X"A7",X"C8",X"11",X"E0",X"FF",X"21",X"E0",X"84",X"3A",X"0E",X"88",X"A7",
		X"28",X"22",X"36",X"02",X"CD",X"AA",X"02",X"21",X"40",X"87",X"CD",X"A8",X"02",X"3A",X"0D",X"88",
		X"A7",X"21",X"40",X"87",X"28",X"03",X"21",X"E0",X"84",X"CB",X"60",X"C8",X"3A",X"06",X"88",X"0F",
		X"D0",X"C3",X"B1",X"02",X"21",X"E0",X"84",X"CD",X"B1",X"02",X"21",X"21",X"85",X"CD",X"B1",X"02",
		X"CD",X"B1",X"02",X"CD",X"B1",X"02",X"18",X"CF",X"36",X"01",X"19",X"36",X"25",X"19",X"36",X"20",
		X"C9",X"3E",X"10",X"77",X"19",X"77",X"19",X"77",X"C9",X"21",X"40",X"88",X"06",X"60",X"AF",X"D7",
		X"21",X"80",X"8A",X"D7",X"D7",X"06",X"37",X"D7",X"C9",X"CD",X"B9",X"02",X"06",X"1D",X"3E",X"20",
		X"90",X"5F",X"16",X"00",X"2A",X"0B",X"88",X"3E",X"10",X"D7",X"19",X"22",X"0B",X"88",X"21",X"09",
		X"88",X"35",X"C9",X"21",X"02",X"84",X"22",X"0B",X"88",X"3E",X"20",X"32",X"09",X"88",X"C9",X"21",
		X"40",X"88",X"DD",X"21",X"80",X"8A",X"11",X"18",X"00",X"06",X"02",X"CD",X"2A",X"03",X"DD",X"21",
		X"90",X"8C",X"06",X"02",X"CD",X"2A",X"03",X"DD",X"21",X"E0",X"8A",X"06",X"12",X"CD",X"43",X"03",
		X"DD",X"21",X"B0",X"8A",X"06",X"02",X"CD",X"2A",X"03",X"21",X"98",X"88",X"35",X"21",X"9C",X"88",
		X"35",X"3A",X"1F",X"88",X"A7",X"C0",X"CD",X"78",X"03",X"C9",X"DD",X"7E",X"06",X"77",X"2C",X"DD",
		X"7E",X"10",X"77",X"2C",X"DD",X"7E",X"04",X"77",X"2C",X"DD",X"7E",X"0F",X"77",X"2C",X"DD",X"19",
		X"10",X"E8",X"C9",X"DD",X"4E",X"05",X"DD",X"7E",X"06",X"CB",X"01",X"17",X"CB",X"01",X"17",X"CB",
		X"01",X"17",X"D6",X"08",X"77",X"2C",X"DD",X"7E",X"10",X"77",X"2C",X"DD",X"7E",X"04",X"DD",X"4E",
		X"03",X"CB",X"01",X"17",X"CB",X"01",X"17",X"CB",X"01",X"17",X"D6",X"08",X"77",X"2C",X"DD",X"7E",
		X"0F",X"77",X"2C",X"DD",X"19",X"10",X"CC",X"C9",X"11",X"40",X"88",X"06",X"18",X"1A",X"ED",X"44",
		X"D6",X"10",X"12",X"1C",X"1A",X"E6",X"C0",X"EE",X"C0",X"4F",X"1A",X"E6",X"0F",X"B1",X"12",X"1C",
		X"1A",X"ED",X"44",X"D6",X"10",X"12",X"1C",X"1C",X"10",X"E3",X"C9",X"3A",X"06",X"88",X"A7",X"C8",
		X"21",X"82",X"84",X"11",X"20",X"00",X"3A",X"80",X"8A",X"3C",X"FE",X"08",X"38",X"02",X"3E",X"08",
		X"4F",X"47",X"36",X"0C",X"19",X"10",X"FB",X"3E",X"08",X"91",X"C8",X"47",X"36",X"10",X"19",X"10",
		X"FB",X"C9",X"21",X"3F",X"86",X"11",X"E0",X"FF",X"3A",X"08",X"89",X"A7",X"C8",X"3D",X"4F",X"28",
		X"0D",X"FE",X"05",X"38",X"02",X"3E",X"05",X"4F",X"47",X"36",X"B0",X"19",X"10",X"FB",X"3E",X"05",
		X"91",X"C8",X"47",X"36",X"10",X"19",X"10",X"FB",X"C9",X"3E",X"1A",X"06",X"0B",X"F5",X"C5",X"CD",
		X"B2",X"05",X"C1",X"F1",X"3C",X"10",X"F6",X"21",X"C7",X"85",X"11",X"20",X"00",X"06",X"0A",X"DD",
		X"21",X"00",X"8A",X"CD",X"29",X"04",X"77",X"19",X"DD",X"23",X"CD",X"29",X"04",X"77",X"19",X"DD",
		X"23",X"CD",X"29",X"04",X"28",X"01",X"77",X"11",X"62",X"FF",X"19",X"11",X"20",X"00",X"DD",X"23",
		X"10",X"E1",X"CD",X"39",X"04",X"CD",X"60",X"04",X"C9",X"DD",X"7E",X"00",X"4F",X"E6",X"0F",X"77",
		X"19",X"79",X"0F",X"0F",X"0F",X"0F",X"E6",X"0F",X"C9",X"DD",X"21",X"C0",X"89",X"21",X"67",X"84",
		X"06",X"0A",X"11",X"20",X"00",X"DD",X"23",X"CD",X"29",X"04",X"77",X"19",X"36",X"51",X"19",X"DD",
		X"23",X"CD",X"29",X"04",X"28",X"01",X"77",X"DD",X"23",X"11",X"82",X"FF",X"19",X"10",X"E3",X"C9",
		X"DD",X"21",X"00",X"8E",X"21",X"67",X"85",X"06",X"0A",X"11",X"E0",X"FF",X"DD",X"7E",X"00",X"A7",
		X"20",X"02",X"3E",X"40",X"77",X"19",X"DD",X"23",X"DD",X"7E",X"00",X"A7",X"20",X"02",X"3E",X"40",
		X"77",X"19",X"DD",X"23",X"DD",X"7E",X"00",X"A7",X"20",X"02",X"3E",X"40",X"77",X"DD",X"23",X"11",
		X"42",X"00",X"19",X"10",X"D4",X"C9",X"4F",X"3A",X"06",X"88",X"0F",X"D0",X"79",X"A7",X"28",X"47",
		X"CD",X"F2",X"04",X"87",X"81",X"4F",X"06",X"00",X"21",X"01",X"05",X"09",X"A7",X"06",X"03",X"1A",
		X"8E",X"27",X"12",X"13",X"23",X"10",X"F8",X"D5",X"3A",X"0D",X"88",X"0F",X"30",X"02",X"3E",X"01",
		X"CD",X"6B",X"05",X"D1",X"1B",X"21",X"AA",X"88",X"06",X"03",X"1A",X"BE",X"D8",X"20",X"05",X"1B",
		X"2B",X"10",X"F7",X"C9",X"CD",X"F2",X"04",X"21",X"A8",X"88",X"06",X"03",X"1A",X"77",X"13",X"23",
		X"10",X"FA",X"3E",X"02",X"C3",X"6B",X"05",X"CD",X"F2",X"04",X"21",X"AB",X"88",X"A7",X"06",X"03",
		X"18",X"BD",X"F5",X"3A",X"0D",X"88",X"11",X"A2",X"88",X"0F",X"30",X"03",X"11",X"A5",X"88",X"F1",
		X"C9",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"07",X"00",X"00",X"05",X"00",X"50",X"04",X"00",
		X"00",X"04",X"00",X"80",X"03",X"00",X"50",X"03",X"00",X"30",X"03",X"00",X"00",X"03",X"00",X"80",
		X"02",X"00",X"50",X"02",X"00",X"30",X"02",X"00",X"00",X"02",X"00",X"80",X"01",X"00",X"50",X"01",
		X"00",X"30",X"01",X"00",X"00",X"01",X"00",X"50",X"00",X"00",X"00",X"01",X"00",X"00",X"01",X"00",
		X"00",X"02",X"00",X"00",X"04",X"00",X"00",X"08",X"00",X"00",X"16",X"00",X"00",X"32",X"00",X"00",
		X"50",X"00",X"F5",X"21",X"A2",X"88",X"A7",X"28",X"09",X"21",X"A5",X"88",X"3D",X"28",X"03",X"21",
		X"A8",X"88",X"36",X"00",X"23",X"36",X"00",X"23",X"36",X"00",X"F1",X"21",X"A4",X"88",X"DD",X"21",
		X"81",X"87",X"A7",X"28",X"11",X"21",X"A7",X"88",X"DD",X"21",X"21",X"85",X"3D",X"28",X"07",X"21",
		X"AA",X"88",X"DD",X"21",X"41",X"86",X"11",X"E0",X"FF",X"06",X"03",X"0E",X"04",X"7E",X"0F",X"0F",
		X"0F",X"0F",X"CD",X"9D",X"05",X"7E",X"CD",X"9D",X"05",X"2B",X"10",X"F1",X"C9",X"E6",X"0F",X"28",
		X"08",X"0E",X"00",X"DD",X"77",X"00",X"DD",X"19",X"C9",X"79",X"A7",X"28",X"F6",X"3E",X"10",X"0D",
		X"18",X"F1",X"87",X"F5",X"21",X"0D",X"7A",X"E6",X"7F",X"5F",X"16",X"00",X"19",X"F1",X"5E",X"23",
		X"56",X"EB",X"5E",X"23",X"56",X"23",X"EB",X"01",X"E0",X"FF",X"38",X"14",X"1A",X"FE",X"2E",X"28",
		X"0B",X"FE",X"3F",X"C8",X"D6",X"30",X"77",X"13",X"09",X"18",X"F1",X"37",X"EB",X"23",X"18",X"E2",
		X"1A",X"FE",X"2E",X"28",X"F6",X"FE",X"3F",X"C8",X"36",X"10",X"13",X"09",X"18",X"F2",X"3E",X"05",
		X"CD",X"B2",X"05",X"3A",X"02",X"88",X"FE",X"63",X"38",X"02",X"3E",X"63",X"CD",X"2A",X"06",X"47",
		X"E6",X"F0",X"28",X"07",X"0F",X"0F",X"0F",X"0F",X"32",X"BF",X"86",X"78",X"E6",X"0F",X"32",X"9F",
		X"86",X"FE",X"02",X"C0",X"11",X"C8",X"64",X"01",X"1F",X"00",X"1A",X"1B",X"80",X"47",X"0D",X"20",
		X"F9",X"FE",X"8C",X"C8",X"21",X"1E",X"45",X"29",X"34",X"C9",X"47",X"E6",X"0F",X"C6",X"00",X"27",
		X"4F",X"78",X"E6",X"F0",X"28",X"0B",X"0F",X"0F",X"0F",X"0F",X"47",X"AF",X"C6",X"16",X"27",X"10",
		X"FB",X"81",X"27",X"C9",X"DD",X"21",X"8A",X"77",X"16",X"00",X"DD",X"7E",X"00",X"FE",X"C8",X"20",
		X"16",X"DD",X"86",X"01",X"30",X"01",X"14",X"DD",X"86",X"02",X"30",X"01",X"14",X"DD",X"86",X"03",
		X"30",X"01",X"14",X"92",X"FE",X"59",X"C8",X"3E",X"01",X"32",X"F8",X"8D",X"C9",X"F5",X"C5",X"D5",
		X"E5",X"08",X"D9",X"F5",X"C5",X"D5",X"E5",X"DD",X"E5",X"FD",X"E5",X"AF",X"32",X"80",X"A1",X"21",
		X"40",X"88",X"DD",X"21",X"10",X"94",X"11",X"10",X"90",X"06",X"04",X"3A",X"0A",X"88",X"FE",X"04",
		X"28",X"04",X"06",X"18",X"18",X"18",X"CD",X"14",X"07",X"21",X"7C",X"88",X"06",X"03",X"CD",X"14",
		X"07",X"21",X"50",X"88",X"06",X"0B",X"CD",X"14",X"07",X"21",X"88",X"88",X"06",X"06",X"CD",X"14",
		X"07",X"32",X"00",X"A0",X"3A",X"15",X"88",X"32",X"16",X"88",X"3A",X"13",X"88",X"32",X"15",X"88",
		X"2A",X"10",X"88",X"22",X"13",X"88",X"21",X"12",X"88",X"3A",X"C0",X"A0",X"2F",X"77",X"2B",X"3A",
		X"A0",X"A0",X"2F",X"77",X"2B",X"3A",X"80",X"A0",X"2F",X"77",X"21",X"3F",X"88",X"35",X"21",X"5F",
		X"8A",X"35",X"CD",X"E8",X"59",X"CD",X"64",X"0E",X"21",X"FA",X"06",X"E5",X"3A",X"05",X"88",X"EF",
		X"2D",X"07",X"99",X"08",X"4E",X"0C",X"9B",X"15",X"53",X"0E",X"3A",X"1F",X"88",X"32",X"87",X"A1",
		X"FD",X"E1",X"DD",X"E1",X"E1",X"D1",X"C1",X"F1",X"D9",X"08",X"E1",X"D1",X"C1",X"3E",X"01",X"32",
		X"80",X"A1",X"F1",X"C9",X"7E",X"DD",X"77",X"01",X"2C",X"7E",X"DD",X"77",X"00",X"2C",X"7E",X"12",
		X"13",X"2C",X"7E",X"12",X"13",X"2C",X"DD",X"23",X"DD",X"23",X"10",X"E8",X"C9",X"06",X"20",X"CD",
		X"CE",X"02",X"C0",X"3A",X"FF",X"8F",X"FE",X"10",X"C2",X"0F",X"02",X"21",X"06",X"88",X"36",X"00",
		X"2B",X"36",X"01",X"AF",X"32",X"0A",X"88",X"01",X"79",X"07",X"CD",X"5D",X"07",X"11",X"04",X"06",
		X"FF",X"11",X"00",X"05",X"FF",X"1E",X"02",X"FF",X"AF",X"32",X"51",X"8E",X"C9",X"21",X"40",X"80",
		X"11",X"20",X"00",X"0A",X"77",X"19",X"7C",X"FE",X"84",X"38",X"F8",X"26",X"80",X"CB",X"F5",X"03",
		X"2C",X"7D",X"E6",X"1F",X"FE",X"1F",X"38",X"EB",X"C9",X"1D",X"03",X"10",X"10",X"17",X"17",X"16",
		X"17",X"17",X"17",X"17",X"17",X"00",X"18",X"18",X"18",X"10",X"10",X"10",X"1B",X"1B",X"1B",X"1B",
		X"1B",X"1B",X"1B",X"1B",X"1B",X"19",X"16",X"16",X"11",X"0D",X"03",X"00",X"00",X"00",X"00",X"00",
		X"00",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",
		X"0A",X"0A",X"0A",X"0A",X"0A",X"00",X"00",X"04",X"00",X"0D",X"03",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"07",X"07",X"00",X"08",X"08",X"08",X"0C",X"0C",X"0C",X"0C",X"0C",X"0E",X"0E",X"0E",X"07",X"07",
		X"07",X"17",X"17",X"17",X"14",X"0E",X"16",X"14",X"00",X"0D",X"03",X"00",X"00",X"0D",X"00",X"00",
		X"07",X"07",X"07",X"07",X"00",X"00",X"00",X"00",X"08",X"08",X"08",X"08",X"0B",X"0B",X"0B",X"0B",
		X"0C",X"0C",X"0C",X"0C",X"00",X"11",X"00",X"04",X"00",X"1D",X"03",X"14",X"11",X"1C",X"1C",X"1C",
		X"1C",X"1C",X"1C",X"1C",X"1C",X"1C",X"1C",X"1C",X"1C",X"1C",X"1C",X"1C",X"1C",X"1C",X"1C",X"1C",
		X"1C",X"1C",X"1C",X"1C",X"1C",X"1F",X"16",X"14",X"11",X"1D",X"03",X"14",X"14",X"00",X"00",X"00",
		X"00",X"00",X"00",X"01",X"01",X"01",X"01",X"01",X"01",X"1B",X"00",X"0C",X"00",X"08",X"00",X"0C",
		X"00",X"19",X"00",X"0E",X"11",X"1F",X"1F",X"10",X"07",X"1D",X"03",X"10",X"10",X"10",X"10",X"10",
		X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",
		X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"11",X"0D",X"03",X"00",X"00",X"07",X"07",X"07",
		X"07",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"0B",X"0B",X"0B",X"0B",X"07",X"00",X"04",X"00",X"1D",X"03",X"12",X"12",X"12",X"12",X"12",
		X"12",X"12",X"12",X"12",X"12",X"12",X"12",X"12",X"12",X"12",X"12",X"12",X"12",X"12",X"12",X"12",
		X"12",X"12",X"12",X"12",X"12",X"12",X"10",X"10",X"11",X"21",X"B5",X"0B",X"E5",X"3A",X"51",X"8E",
		X"EF",X"B3",X"08",X"E9",X"08",X"2C",X"09",X"86",X"09",X"9C",X"09",X"C8",X"0A",X"32",X"0B",X"42",
		X"74",X"EA",X"76",X"AF",X"32",X"28",X"A0",X"32",X"19",X"88",X"CD",X"E3",X"02",X"21",X"51",X"8E",
		X"34",X"01",X"D5",X"64",X"2E",X"00",X"65",X"0A",X"FE",X"96",X"28",X"08",X"84",X"30",X"01",X"2C",
		X"67",X"0B",X"18",X"F3",X"95",X"FE",X"8F",X"28",X"05",X"3E",X"01",X"32",X"FB",X"89",X"AF",X"32",
		X"06",X"88",X"CD",X"B9",X"02",X"CD",X"0D",X"1D",X"C9",X"06",X"1D",X"CD",X"CE",X"02",X"C0",X"CD",
		X"E3",X"02",X"21",X"59",X"08",X"06",X"1F",X"7E",X"23",X"86",X"10",X"FC",X"FE",X"63",X"20",X"F2",
		X"01",X"59",X"08",X"CD",X"5D",X"07",X"21",X"31",X"08",X"06",X"08",X"7E",X"23",X"86",X"10",X"FC",
		X"FE",X"AA",X"20",X"DE",X"CD",X"54",X"0E",X"11",X"11",X"06",X"FF",X"1E",X"0B",X"FF",X"21",X"51",
		X"8E",X"36",X"07",X"C9",X"58",X"40",X"38",X"06",X"88",X"40",X"38",X"0B",X"06",X"19",X"CD",X"CE",
		X"02",X"C0",X"CD",X"E3",X"02",X"21",X"51",X"8E",X"34",X"CD",X"B9",X"02",X"21",X"F5",X"07",X"3E",
		X"11",X"BE",X"20",X"FD",X"DD",X"21",X"38",X"08",X"06",X"07",X"21",X"76",X"09",X"78",X"CD",X"45",
		X"0C",X"3E",X"1C",X"83",X"5F",X"30",X"01",X"14",X"1A",X"4F",X"DD",X"7E",X"00",X"B9",X"20",X"16",
		X"DD",X"2B",X"10",X"E6",X"01",X"D9",X"07",X"CD",X"5D",X"07",X"11",X"8B",X"06",X"FF",X"1E",X"8E",
		X"FF",X"11",X"00",X"02",X"FF",X"C9",X"79",X"07",X"99",X"07",X"B9",X"07",X"D9",X"07",X"F9",X"07",
		X"19",X"08",X"39",X"08",X"59",X"08",X"21",X"50",X"8E",X"35",X"C0",X"CD",X"B9",X"02",X"CD",X"E3",
		X"02",X"21",X"51",X"8E",X"34",X"21",X"26",X"0B",X"22",X"48",X"8F",X"C9",X"06",X"19",X"CD",X"CE",
		X"02",X"C0",X"16",X"0D",X"21",X"65",X"0A",X"01",X"C9",X"07",X"0A",X"96",X"20",X"FC",X"03",X"23",
		X"15",X"20",X"F7",X"01",X"B9",X"07",X"CD",X"5D",X"07",X"11",X"0D",X"06",X"FF",X"21",X"70",X"8B",
		X"AF",X"47",X"D7",X"21",X"76",X"0A",X"11",X"7E",X"0A",X"DD",X"21",X"70",X"8B",X"CD",X"0C",X"0A",
		X"01",X"18",X"00",X"DD",X"09",X"1A",X"3C",X"20",X"F4",X"CD",X"52",X"0A",X"CD",X"25",X"0A",X"21",
		X"87",X"0A",X"22",X"54",X"8E",X"21",X"48",X"86",X"22",X"56",X"8E",X"21",X"50",X"8E",X"36",X"32",
		X"2C",X"34",X"2C",X"36",X"0D",X"2C",X"36",X"05",X"DD",X"21",X"70",X"8B",X"06",X"04",X"11",X"18",
		X"00",X"CD",X"06",X"40",X"DD",X"19",X"10",X"F9",X"CD",X"EF",X"02",X"C9",X"1A",X"DD",X"77",X"06",
		X"13",X"1A",X"13",X"DD",X"77",X"04",X"7E",X"DD",X"77",X"0C",X"23",X"7E",X"DD",X"77",X"0D",X"DD",
		X"36",X"0E",X"00",X"23",X"C9",X"21",X"41",X"8D",X"36",X"0A",X"2D",X"7E",X"34",X"E6",X"03",X"21",
		X"F6",X"26",X"CD",X"45",X"0C",X"D5",X"21",X"6A",X"86",X"CD",X"40",X"0A",X"D1",X"21",X"AA",X"86",
		X"01",X"20",X"00",X"1A",X"77",X"2C",X"13",X"1A",X"77",X"09",X"13",X"1A",X"77",X"2D",X"13",X"1A",
		X"77",X"C9",X"21",X"AA",X"82",X"11",X"72",X"0A",X"CD",X"40",X"0A",X"21",X"6A",X"82",X"11",X"72",
		X"0A",X"CD",X"40",X"0A",X"C9",X"0C",X"0C",X"0E",X"0E",X"0E",X"07",X"07",X"07",X"17",X"17",X"17",
		X"14",X"0E",X"00",X"00",X"00",X"00",X"5D",X"2D",X"EF",X"68",X"38",X"38",X"12",X"42",X"0A",X"08",
		X"0A",X"0E",X"0A",X"13",X"0A",X"16",X"FF",X"10",X"40",X"40",X"40",X"10",X"10",X"20",X"1F",X"1F",
		X"29",X"11",X"1E",X"10",X"10",X"40",X"40",X"40",X"10",X"10",X"12",X"25",X"25",X"29",X"11",X"1E",
		X"10",X"10",X"40",X"40",X"40",X"10",X"10",X"1D",X"11",X"1D",X"11",X"10",X"10",X"10",X"10",X"40",
		X"40",X"40",X"10",X"10",X"27",X"1F",X"1C",X"16",X"10",X"10",X"10",X"10",X"40",X"40",X"40",X"10",
		X"10",X"12",X"1F",X"23",X"23",X"10",X"10",X"10",X"21",X"41",X"8D",X"35",X"20",X"03",X"CD",X"28",
		X"0A",X"CD",X"F8",X"09",X"21",X"50",X"8E",X"35",X"C0",X"36",X"02",X"2A",X"54",X"8E",X"7E",X"23",
		X"22",X"54",X"8E",X"2A",X"56",X"8E",X"77",X"11",X"E0",X"FF",X"19",X"22",X"56",X"8E",X"21",X"52",
		X"8E",X"35",X"C0",X"36",X"0D",X"21",X"50",X"8E",X"36",X"14",X"2C",X"34",X"2A",X"56",X"8E",X"11",
		X"00",X"00",X"06",X"0E",X"7E",X"83",X"5F",X"30",X"01",X"14",X"3E",X"20",X"85",X"6F",X"30",X"01",
		X"24",X"10",X"F1",X"2A",X"48",X"8F",X"7E",X"BB",X"C2",X"42",X"74",X"23",X"7E",X"BA",X"C2",X"EA",
		X"76",X"23",X"22",X"48",X"8F",X"C9",X"C6",X"01",X"C4",X"01",X"8C",X"01",X"A8",X"01",X"A7",X"01",
		X"BC",X"1C",X"21",X"BC",X"82",X"11",X"E0",X"FF",X"06",X"0A",X"7E",X"19",X"BE",X"C2",X"B3",X"08",
		X"10",X"F8",X"21",X"41",X"8D",X"35",X"20",X"03",X"CD",X"28",X"0A",X"CD",X"F8",X"09",X"21",X"50",
		X"8E",X"35",X"C0",X"36",X"01",X"2C",X"35",X"3A",X"53",X"8E",X"3D",X"21",X"AB",X"0B",X"CD",X"45",
		X"0C",X"ED",X"53",X"56",X"8E",X"21",X"53",X"8E",X"35",X"C0",X"21",X"50",X"8E",X"36",X"96",X"2C",
		X"AF",X"77",X"21",X"62",X"84",X"57",X"5F",X"0E",X"0E",X"06",X"1D",X"7B",X"86",X"30",X"01",X"14",
		X"5F",X"23",X"10",X"F7",X"7D",X"C6",X"03",X"6F",X"30",X"01",X"24",X"0D",X"20",X"EB",X"2A",X"48",
		X"8F",X"7B",X"BE",X"C2",X"B3",X"08",X"23",X"7E",X"BA",X"C2",X"E9",X"08",X"AF",X"32",X"48",X"8F",
		X"32",X"49",X"8F",X"3E",X"03",X"32",X"05",X"88",X"C3",X"00",X"0E",X"59",X"86",X"56",X"86",X"53",
		X"86",X"4E",X"86",X"4B",X"86",X"3A",X"06",X"88",X"A7",X"20",X"41",X"3A",X"05",X"88",X"3D",X"20",
		X"3B",X"3A",X"51",X"8E",X"FE",X"03",X"28",X"08",X"FE",X"05",X"28",X"04",X"FE",X"08",X"20",X"2C",
		X"11",X"E0",X"FF",X"21",X"FE",X"8E",X"34",X"21",X"BC",X"86",X"01",X"C2",X"20",X"0A",X"96",X"20",
		X"16",X"19",X"03",X"0A",X"3C",X"20",X"F6",X"11",X"C0",X"FB",X"19",X"EB",X"21",X"CB",X"20",X"3A",
		X"51",X"8E",X"E7",X"EB",X"BE",X"28",X"05",X"3E",X"01",X"32",X"E5",X"89",X"3A",X"2C",X"88",X"FE",
		X"0F",X"20",X"19",X"3A",X"10",X"88",X"CB",X"5F",X"28",X"09",X"CD",X"CF",X"0E",X"21",X"00",X"00",
		X"C3",X"AB",X"0D",X"CB",X"67",X"C8",X"CD",X"CF",X"0E",X"C3",X"A8",X"0D",X"3A",X"02",X"88",X"A7",
		X"C8",X"21",X"05",X"88",X"34",X"AF",X"32",X"0A",X"88",X"C9",X"3A",X"80",X"A0",X"CB",X"5F",X"C0",
		X"3E",X"09",X"32",X"51",X"8E",X"21",X"00",X"84",X"1E",X"10",X"01",X"FF",X"03",X"73",X"23",X"0B",
		X"78",X"B1",X"20",X"F9",X"C9",X"87",X"16",X"00",X"5F",X"19",X"5E",X"23",X"56",X"C9",X"21",X"78",
		X"0D",X"E5",X"3A",X"0A",X"88",X"EF",X"5C",X"0C",X"77",X"0C",X"61",X"0D",X"AF",X"32",X"19",X"88",
		X"32",X"28",X"A0",X"32",X"06",X"88",X"21",X"42",X"84",X"22",X"0B",X"88",X"21",X"09",X"88",X"36",
		X"0F",X"23",X"34",X"CD",X"B9",X"02",X"C9",X"2A",X"0B",X"88",X"06",X"1D",X"3E",X"10",X"D7",X"11",
		X"03",X"00",X"19",X"06",X"1D",X"D7",X"19",X"22",X"0B",X"88",X"21",X"09",X"88",X"35",X"C0",X"2C",
		X"34",X"21",X"79",X"07",X"01",X"00",X"00",X"7E",X"23",X"86",X"30",X"01",X"0C",X"10",X"F9",X"FE",
		X"C1",X"20",X"F5",X"79",X"FE",X"0C",X"20",X"F0",X"01",X"79",X"07",X"CD",X"5D",X"07",X"32",X"0D",
		X"88",X"CD",X"54",X"0E",X"CD",X"F8",X"0C",X"11",X"01",X"06",X"FF",X"1E",X"11",X"FF",X"1E",X"16",
		X"FF",X"1C",X"3A",X"00",X"88",X"E6",X"01",X"28",X"02",X"1E",X"28",X"FF",X"1E",X"2A",X"3A",X"00",
		X"88",X"E6",X"01",X"28",X"01",X"1D",X"FF",X"CD",X"4E",X"0F",X"21",X"26",X"0B",X"11",X"00",X"00",
		X"06",X"20",X"7E",X"83",X"5F",X"30",X"01",X"14",X"23",X"10",X"F7",X"7B",X"FE",X"D3",X"00",X"00",
		X"00",X"3E",X"0B",X"BA",X"00",X"00",X"00",X"C9",X"21",X"2F",X"0D",X"DD",X"21",X"A7",X"86",X"11",
		X"E0",X"FF",X"06",X"0C",X"7E",X"DD",X"77",X"00",X"23",X"DD",X"19",X"10",X"F7",X"7E",X"FE",X"FF",
		X"28",X"0F",X"FE",X"EE",X"C8",X"11",X"81",X"01",X"DD",X"19",X"11",X"E0",X"FF",X"06",X"0C",X"18",
		X"E3",X"21",X"48",X"0D",X"DD",X"21",X"A7",X"82",X"11",X"E0",X"FF",X"06",X"0C",X"18",X"D5",X"0C",
		X"0C",X"0C",X"0C",X"0C",X"0C",X"0E",X"0E",X"0C",X"0C",X"A4",X"A5",X"0D",X"0C",X"0C",X"0C",X"0C",
		X"0C",X"0F",X"0F",X"3B",X"3B",X"A5",X"A4",X"FF",X"00",X"80",X"03",X"83",X"0D",X"8D",X"00",X"80",
		X"05",X"85",X"00",X"C0",X"00",X"C0",X"43",X"C3",X"4D",X"CD",X"00",X"80",X"02",X"82",X"00",X"C0",
		X"EE",X"3A",X"02",X"88",X"A7",X"C8",X"3D",X"11",X"18",X"06",X"28",X"01",X"1C",X"FF",X"11",X"00",
		X"03",X"FF",X"3E",X"02",X"32",X"05",X"88",X"C9",X"3A",X"10",X"88",X"CB",X"5F",X"C2",X"E4",X"0D",
		X"CB",X"67",X"C8",X"3A",X"02",X"88",X"FE",X"02",X"D8",X"D6",X"02",X"32",X"02",X"88",X"21",X"6B",
		X"77",X"06",X"14",X"58",X"53",X"7E",X"83",X"5F",X"30",X"01",X"14",X"23",X"10",X"F7",X"7B",X"82",
		X"E6",X"AB",X"28",X"04",X"21",X"EA",X"89",X"34",X"21",X"00",X"01",X"22",X"0D",X"88",X"CD",X"54",
		X"0E",X"AF",X"32",X"0A",X"88",X"3E",X"03",X"32",X"05",X"88",X"3E",X"01",X"32",X"06",X"88",X"32",
		X"1F",X"88",X"11",X"04",X"06",X"FF",X"CD",X"00",X"0E",X"21",X"21",X"8D",X"36",X"00",X"2C",X"36",
		X"20",X"11",X"00",X"04",X"FF",X"3A",X"0E",X"88",X"0F",X"D0",X"1C",X"FF",X"AF",X"21",X"1F",X"8E",
		X"06",X"0C",X"D7",X"C9",X"3A",X"02",X"88",X"A7",X"28",X"0A",X"3D",X"32",X"02",X"88",X"21",X"00",
		X"00",X"C3",X"AB",X"0D",X"3A",X"0A",X"88",X"FE",X"0E",X"C8",X"3E",X"01",X"32",X"05",X"88",X"C9",
		X"21",X"00",X"89",X"AF",X"32",X"0A",X"88",X"32",X"E1",X"89",X"32",X"E2",X"89",X"32",X"E3",X"89",
		X"32",X"5B",X"8F",X"06",X"BF",X"D7",X"3A",X"07",X"88",X"32",X"48",X"89",X"32",X"88",X"89",X"3E",
		X"20",X"32",X"41",X"89",X"32",X"81",X"89",X"3A",X"20",X"88",X"32",X"40",X"89",X"32",X"80",X"89",
		X"CD",X"E3",X"02",X"3A",X"06",X"88",X"A7",X"C8",X"AF",X"32",X"3F",X"8F",X"32",X"30",X"8F",X"32",
		X"0E",X"8F",X"32",X"0F",X"8F",X"C9",X"11",X"04",X"00",X"06",X"06",X"3E",X"FB",X"A6",X"77",X"19",
		X"10",X"F9",X"C9",X"C9",X"11",X"01",X"07",X"FF",X"3A",X"2C",X"88",X"FE",X"0F",X"20",X"04",X"11",
		X"06",X"06",X"FF",X"C9",X"11",X"41",X"8A",X"1A",X"6F",X"26",X"8A",X"7E",X"FE",X"FF",X"C8",X"47",
		X"3A",X"21",X"88",X"E6",X"01",X"20",X"06",X"3A",X"06",X"88",X"A7",X"28",X"04",X"78",X"CD",X"8F",
		X"0E",X"36",X"FF",X"7D",X"FE",X"5E",X"28",X"03",X"3C",X"12",X"C9",X"3E",X"43",X"12",X"C9",X"32",
		X"00",X"A1",X"3E",X"01",X"32",X"81",X"A1",X"00",X"00",X"00",X"00",X"00",X"00",X"3D",X"32",X"81",
		X"A1",X"C9",X"32",X"20",X"8D",X"3A",X"06",X"88",X"A7",X"20",X"05",X"3A",X"50",X"8F",X"A7",X"C8",
		X"3A",X"20",X"8D",X"C5",X"D5",X"E5",X"47",X"11",X"40",X"8A",X"1A",X"6F",X"26",X"8A",X"70",X"7D",
		X"FE",X"5E",X"28",X"04",X"3C",X"12",X"18",X"03",X"3E",X"43",X"12",X"E1",X"D1",X"C1",X"C9",X"AF",
		X"18",X"E1",X"3E",X"01",X"18",X"CC",X"3E",X"02",X"18",X"D9",X"3E",X"82",X"CD",X"B3",X"0E",X"3E",
		X"03",X"18",X"D0",X"3A",X"24",X"8F",X"A7",X"C0",X"3A",X"32",X"8D",X"A7",X"C0",X"3E",X"04",X"18",
		X"B1",X"3E",X"05",X"18",X"BE",X"3E",X"06",X"18",X"A9",X"3E",X"07",X"18",X"A5",X"3E",X"08",X"18",
		X"A1",X"3E",X"09",X"18",X"AE",X"3E",X"0A",X"18",X"99",X"3E",X"0B",X"18",X"82",X"3E",X"0B",X"18",
		X"91",X"3E",X"0C",X"18",X"8D",X"3E",X"0D",X"18",X"89",X"3E",X"0E",X"18",X"85",X"3E",X"0F",X"18",
		X"81",X"3E",X"95",X"CD",X"A2",X"0E",X"3E",X"10",X"C3",X"A2",X"0E",X"3E",X"11",X"C3",X"A2",X"0E",
		X"3E",X"95",X"CD",X"A2",X"0E",X"3E",X"03",X"CD",X"A2",X"0E",X"3E",X"11",X"C3",X"A2",X"0E",X"3E",
		X"12",X"C3",X"A2",X"0E",X"3E",X"13",X"C3",X"A2",X"0E",X"3E",X"14",X"C3",X"A2",X"0E",X"3E",X"82",
		X"CD",X"B3",X"0E",X"3E",X"95",X"C3",X"B3",X"0E",X"3E",X"96",X"CD",X"A2",X"0E",X"3E",X"97",X"CD",
		X"A2",X"0E",X"3E",X"18",X"CD",X"B3",X"0E",X"3E",X"15",X"C3",X"B3",X"0E",X"3E",X"19",X"CD",X"B3",
		X"0E",X"3E",X"15",X"C3",X"B3",X"0E",X"3A",X"68",X"8D",X"B7",X"C0",X"3A",X"07",X"89",X"E6",X"01",
		X"C6",X"1A",X"CD",X"A2",X"0E",X"C3",X"C3",X"0F",X"3E",X"82",X"CD",X"A2",X"0E",X"3E",X"1C",X"C3",
		X"C3",X"0F",X"3E",X"1D",X"C3",X"C3",X"0F",X"3A",X"07",X"89",X"0F",X"E6",X"03",X"C6",X"1E",X"C3",
		X"C3",X"0F",X"3A",X"07",X"89",X"0F",X"E6",X"03",X"C6",X"22",X"C3",X"C3",X"0F",X"3E",X"26",X"C3",
		X"C3",X"0F",X"3E",X"27",X"CD",X"B3",X"0E",X"3E",X"15",X"C3",X"B3",X"0E",X"3E",X"28",X"C3",X"C3",
		X"0F",X"3E",X"29",X"CD",X"A2",X"0E",X"3E",X"15",X"CD",X"A2",X"0E",X"3E",X"16",X"CD",X"A2",X"0E",
		X"3E",X"17",X"C3",X"A2",X"0E",X"3A",X"5C",X"8F",X"E6",X"07",X"FE",X"02",X"38",X"04",X"21",X"35",
		X"10",X"E5",X"EF",X"EF",X"0F",X"16",X"10",X"90",X"10",X"A2",X"10",X"3C",X"11",X"4F",X"11",X"3E",
		X"0F",X"21",X"01",X"89",X"77",X"2E",X"07",X"CB",X"56",X"28",X"03",X"CD",X"F1",X"50",X"3E",X"01",
		X"32",X"61",X"8F",X"32",X"3F",X"8F",X"32",X"5C",X"8F",X"CD",X"BC",X"0F",X"21",X"38",X"8A",X"7E",
		X"23",X"B7",X"C8",X"32",X"5C",X"8F",X"CD",X"83",X"15",X"CD",X"42",X"10",X"CD",X"7D",X"10",X"CD",
		X"D4",X"20",X"CD",X"1B",X"51",X"CD",X"19",X"12",X"CD",X"BD",X"40",X"CD",X"EF",X"02",X"CD",X"E4",
		X"5A",X"CD",X"64",X"0E",X"C9",X"CD",X"57",X"21",X"CD",X"19",X"12",X"CD",X"BD",X"40",X"CD",X"EF",
		X"02",X"C9",X"3E",X"01",X"32",X"3F",X"8F",X"DD",X"21",X"80",X"8A",X"FD",X"21",X"90",X"8C",X"DD",
		X"7E",X"02",X"A7",X"20",X"23",X"3A",X"24",X"8F",X"21",X"57",X"8F",X"B6",X"20",X"1A",X"3A",X"1F",
		X"88",X"A7",X"3A",X"A0",X"A0",X"20",X"03",X"3A",X"C0",X"A0",X"2F",X"DD",X"77",X"07",X"DD",X"7E",
		X"1E",X"A7",X"C0",X"DD",X"CB",X"07",X"A6",X"C9",X"DD",X"36",X"07",X"00",X"C9",X"3A",X"01",X"89",
		X"A7",X"C0",X"21",X"5C",X"8F",X"34",X"11",X"35",X"06",X"FF",X"3E",X"40",X"32",X"62",X"8F",X"C9",
		X"21",X"62",X"8F",X"7E",X"A7",X"28",X"02",X"35",X"C9",X"21",X"5C",X"8F",X"34",X"11",X"34",X"06",
		X"FF",X"C9",X"3A",X"5D",X"8F",X"FE",X"0A",X"38",X"04",X"47",X"CD",X"31",X"11",X"21",X"50",X"86",
		X"CD",X"19",X"11",X"3A",X"5D",X"8F",X"A7",X"28",X"26",X"FE",X"0C",X"30",X"22",X"D6",X"07",X"06",
		X"05",X"28",X"0D",X"30",X"06",X"04",X"3C",X"20",X"FC",X"18",X"05",X"05",X"3D",X"20",X"FC",X"78",
		X"78",X"32",X"62",X"8F",X"CB",X"20",X"CD",X"31",X"11",X"21",X"D0",X"85",X"CD",X"19",X"11",X"3A",
		X"5E",X"8F",X"FE",X"0A",X"38",X"04",X"47",X"CD",X"31",X"11",X"21",X"52",X"86",X"CD",X"19",X"11",
		X"21",X"60",X"8F",X"7E",X"A7",X"28",X"1A",X"47",X"2E",X"62",X"86",X"77",X"CB",X"20",X"CD",X"31",
		X"11",X"5F",X"79",X"A7",X"28",X"04",X"79",X"32",X"F2",X"85",X"21",X"D2",X"85",X"7B",X"CD",X"19",
		X"11",X"21",X"5C",X"8F",X"34",X"CD",X"44",X"0F",X"C9",X"01",X"E0",X"FF",X"5F",X"CB",X"3F",X"CB",
		X"3F",X"CB",X"3F",X"CB",X"3F",X"A7",X"20",X"02",X"3E",X"10",X"77",X"09",X"7B",X"E6",X"0F",X"77",
		X"C9",X"AF",X"4F",X"C6",X"01",X"27",X"30",X"01",X"0C",X"10",X"F8",X"C9",X"21",X"62",X"8F",X"7E",
		X"A7",X"28",X"06",X"35",X"11",X"15",X"03",X"FF",X"C9",X"36",X"80",X"2E",X"5C",X"34",X"C9",X"21",
		X"62",X"8F",X"7E",X"A7",X"28",X"02",X"35",X"C9",X"AF",X"2E",X"5B",X"06",X"09",X"D7",X"CD",X"CF",
		X"0E",X"3E",X"06",X"32",X"0A",X"88",X"21",X"3C",X"8A",X"3A",X"2B",X"88",X"86",X"A7",X"C8",X"18",
		X"1C",X"21",X"07",X"8D",X"7E",X"A7",X"28",X"02",X"35",X"C9",X"3A",X"01",X"89",X"2E",X"40",X"96",
		X"C8",X"D8",X"4F",X"7E",X"FE",X"06",X"D0",X"DD",X"21",X"E0",X"8A",X"06",X"06",X"1E",X"1D",X"CD",
		X"9A",X"11",X"11",X"18",X"00",X"DD",X"19",X"10",X"F4",X"C9",X"DD",X"7E",X"00",X"DD",X"B6",X"01",
		X"0F",X"D8",X"41",X"DD",X"36",X"00",X"01",X"DD",X"36",X"02",X"03",X"DD",X"73",X"04",X"AF",X"DD",
		X"77",X"03",X"DD",X"77",X"05",X"DD",X"77",X"06",X"DD",X"77",X"08",X"DD",X"36",X"07",X"01",X"DD",
		X"77",X"0B",X"21",X"09",X"12",X"3A",X"07",X"89",X"E6",X"3F",X"CB",X"3F",X"CB",X"3F",X"FE",X"10",
		X"E7",X"DD",X"77",X"09",X"ED",X"44",X"DD",X"77",X"0A",X"11",X"29",X"38",X"CD",X"1E",X"38",X"21",
		X"F9",X"11",X"3A",X"07",X"89",X"E6",X"3F",X"CB",X"2F",X"CB",X"2F",X"E7",X"32",X"07",X"8D",X"21",
		X"5F",X"8F",X"34",X"21",X"40",X"8D",X"34",X"F1",X"C9",X"50",X"4C",X"48",X"44",X"40",X"3C",X"38",
		X"30",X"2E",X"2C",X"2A",X"28",X"26",X"24",X"24",X"22",X"14",X"14",X"16",X"16",X"18",X"18",X"1A",
		X"1A",X"1B",X"1B",X"1C",X"1C",X"1D",X"1D",X"1E",X"1E",X"DD",X"21",X"E0",X"8A",X"11",X"18",X"00",
		X"06",X"0E",X"D9",X"CD",X"2C",X"12",X"D9",X"DD",X"19",X"10",X"F7",X"C9",X"DD",X"7E",X"00",X"DD",
		X"B6",X"01",X"0F",X"D0",X"DD",X"7E",X"02",X"E6",X"1F",X"FE",X"11",X"D0",X"EF",X"5F",X"12",X"70",
		X"12",X"36",X"35",X"AF",X"12",X"65",X"38",X"96",X"14",X"E3",X"3B",X"92",X"3C",X"DC",X"14",X"18",
		X"15",X"4D",X"15",X"69",X"3E",X"9C",X"3E",X"5C",X"3F",X"72",X"3F",X"7C",X"3F",X"E9",X"3F",X"DD",
		X"35",X"11",X"C0",X"DD",X"34",X"02",X"11",X"38",X"38",X"DD",X"36",X"08",X"01",X"C3",X"1E",X"38",
		X"CD",X"06",X"40",X"DD",X"7E",X"0A",X"ED",X"44",X"47",X"DD",X"7E",X"05",X"B8",X"30",X"03",X"DD",
		X"35",X"06",X"DD",X"86",X"0A",X"DD",X"77",X"05",X"DD",X"7E",X"06",X"A7",X"C0",X"CD",X"53",X"35",
		X"21",X"40",X"8D",X"35",X"21",X"01",X"89",X"7E",X"4F",X"A7",X"28",X"01",X"35",X"3A",X"0A",X"88",
		X"FE",X"04",X"20",X"02",X"2C",X"34",X"79",X"3D",X"FE",X"0A",X"D0",X"32",X"43",X"87",X"C9",X"CD",
		X"06",X"40",X"DD",X"7E",X"08",X"A7",X"C2",X"FE",X"13",X"DD",X"7E",X"05",X"DD",X"86",X"09",X"30",
		X"03",X"DD",X"34",X"06",X"DD",X"77",X"05",X"47",X"3A",X"01",X"89",X"FE",X"03",X"DA",X"99",X"13",
		X"21",X"FB",X"12",X"3A",X"07",X"89",X"E6",X"1F",X"CB",X"3F",X"CB",X"3F",X"CD",X"45",X"0C",X"EB",
		X"3A",X"41",X"8D",X"E6",X"0F",X"E7",X"4F",X"DD",X"7E",X"06",X"B9",X"CA",X"83",X"13",X"FE",X"14",
		X"D8",X"DD",X"36",X"08",X"01",X"11",X"38",X"38",X"C3",X"1E",X"38",X"0B",X"13",X"1A",X"13",X"29",
		X"13",X"38",X"13",X"47",X"13",X"56",X"13",X"65",X"13",X"74",X"13",X"11",X"0D",X"09",X"0D",X"09",
		X"12",X"0E",X"0B",X"09",X"0D",X"09",X"09",X"11",X"0D",X"09",X"0D",X"09",X"11",X"0D",X"09",X"09",
		X"12",X"10",X"09",X"0D",X"09",X"11",X"0D",X"09",X"09",X"11",X"0D",X"11",X"0D",X"09",X"11",X"0F",
		X"0D",X"09",X"12",X"0D",X"10",X"09",X"0D",X"09",X"09",X"09",X"09",X"11",X"0C",X"08",X"0D",X"09",
		X"11",X"0E",X"0B",X"08",X"11",X"0D",X"09",X"11",X"0D",X"09",X"0D",X"11",X"0D",X"09",X"0D",X"11",
		X"0D",X"09",X"0D",X"11",X"0D",X"09",X"11",X"0D",X"09",X"09",X"11",X"0D",X"0D",X"09",X"12",X"11",
		X"0D",X"09",X"11",X"0D",X"09",X"0D",X"09",X"0B",X"08",X"11",X"12",X"0D",X"11",X"0D",X"10",X"09",
		X"10",X"11",X"0D",X"09",X"11",X"0D",X"0B",X"09",X"12",X"10",X"0D",X"0C",X"09",X"0B",X"10",X"0C",
		X"11",X"0D",X"18",X"78",X"FE",X"20",X"D0",X"18",X"33",X"DD",X"CB",X"08",X"46",X"C8",X"C3",X"1C",
		X"14",X"DD",X"CB",X"08",X"46",X"C0",X"C3",X"D0",X"12",X"DD",X"7E",X"06",X"FE",X"07",X"38",X"E9",
		X"FE",X"14",X"30",X"ED",X"21",X"6B",X"8D",X"7E",X"A7",X"28",X"02",X"35",X"C9",X"78",X"FE",X"80",
		X"D0",X"EB",X"21",X"D3",X"13",X"3A",X"07",X"89",X"E6",X"07",X"E7",X"12",X"FD",X"21",X"70",X"8B",
		X"11",X"18",X"00",X"06",X"05",X"FD",X"7E",X"00",X"FD",X"B6",X"01",X"0F",X"30",X"0D",X"FD",X"19",
		X"10",X"F3",X"C9",X"28",X"28",X"20",X"20",X"18",X"18",X"10",X"10",X"21",X"41",X"8D",X"34",X"20",
		X"01",X"34",X"4E",X"DD",X"71",X"14",X"21",X"88",X"39",X"DD",X"75",X"0C",X"DD",X"74",X"0D",X"DD",
		X"36",X"0E",X"00",X"DD",X"36",X"11",X"28",X"DD",X"36",X"02",X"04",X"C3",X"2C",X"14",X"DD",X"7E",
		X"0A",X"ED",X"44",X"47",X"DD",X"7E",X"05",X"B8",X"30",X"03",X"DD",X"35",X"06",X"DD",X"86",X"0A",
		X"DD",X"77",X"05",X"47",X"3A",X"01",X"89",X"FE",X"03",X"DA",X"99",X"13",X"DD",X"7E",X"06",X"FE",
		X"02",X"D0",X"DD",X"36",X"08",X"00",X"11",X"29",X"38",X"C3",X"1E",X"38",X"FD",X"36",X"00",X"01",
		X"FD",X"36",X"02",X"04",X"FD",X"71",X"14",X"AF",X"FD",X"77",X"07",X"FD",X"77",X"0E",X"DD",X"7E",
		X"05",X"C6",X"80",X"FD",X"77",X"05",X"DD",X"7E",X"03",X"C6",X"80",X"FD",X"77",X"03",X"DD",X"7E",
		X"04",X"D6",X"01",X"FD",X"77",X"04",X"DD",X"7E",X"06",X"C6",X"01",X"FD",X"77",X"06",X"3A",X"00",
		X"89",X"FE",X"08",X"38",X"02",X"3E",X"07",X"21",X"8E",X"14",X"E7",X"3A",X"07",X"89",X"E6",X"01",
		X"7E",X"28",X"02",X"ED",X"44",X"FD",X"77",X"0A",X"DD",X"77",X"0A",X"11",X"CB",X"38",X"FD",X"77",
		X"0B",X"FD",X"73",X"0C",X"FD",X"72",X"0D",X"FD",X"36",X"11",X"28",X"C3",X"E3",X"0E",X"10",X"11",
		X"12",X"13",X"14",X"15",X"16",X"17",X"CD",X"06",X"40",X"DD",X"7E",X"0A",X"ED",X"44",X"47",X"DD",
		X"7E",X"03",X"B8",X"30",X"03",X"DD",X"35",X"04",X"DD",X"86",X"0A",X"DD",X"77",X"03",X"DD",X"46",
		X"04",X"DD",X"7E",X"07",X"A7",X"28",X"12",X"78",X"FE",X"04",X"38",X"04",X"DD",X"7E",X"06",X"C9",
		X"DD",X"36",X"02",X"00",X"DD",X"36",X"11",X"20",X"C9",X"78",X"FE",X"02",X"D0",X"11",X"D1",X"3B",
		X"CD",X"1E",X"38",X"DD",X"36",X"02",X"02",X"DD",X"36",X"11",X"28",X"C9",X"06",X"01",X"DD",X"4E",
		X"17",X"3A",X"45",X"8D",X"A7",X"28",X"21",X"DD",X"4E",X"12",X"0C",X"28",X"1B",X"FE",X"05",X"38",
		X"02",X"3E",X"04",X"47",X"05",X"48",X"28",X"06",X"3E",X"01",X"CB",X"27",X"10",X"FC",X"21",X"60",
		X"8F",X"86",X"77",X"2E",X"5E",X"34",X"06",X"38",X"DD",X"70",X"11",X"79",X"21",X"57",X"15",X"CD",
		X"45",X"0C",X"CD",X"1E",X"38",X"DD",X"34",X"02",X"CD",X"06",X"40",X"DD",X"35",X"11",X"C0",X"3A",
		X"60",X"8F",X"CB",X"27",X"47",X"A7",X"28",X"12",X"CD",X"31",X"11",X"5F",X"79",X"A7",X"28",X"03",
		X"32",X"E9",X"85",X"21",X"C9",X"85",X"7B",X"CD",X"19",X"11",X"DD",X"7E",X"16",X"FE",X"07",X"CA",
		X"99",X"3D",X"3C",X"DD",X"77",X"13",X"DD",X"36",X"11",X"01",X"DD",X"34",X"02",X"CD",X"06",X"40",
		X"DD",X"35",X"11",X"C0",X"C3",X"53",X"35",X"5F",X"15",X"68",X"15",X"71",X"15",X"7A",X"15",X"80",
		X"01",X"05",X"40",X"1D",X"05",X"42",X"37",X"28",X"80",X"01",X"05",X"40",X"1D",X"05",X"43",X"39",
		X"28",X"80",X"01",X"04",X"40",X"1D",X"04",X"42",X"39",X"28",X"80",X"01",X"03",X"40",X"1D",X"03",
		X"4F",X"3A",X"38",X"21",X"4D",X"8F",X"34",X"7E",X"47",X"E6",X"0F",X"C0",X"CB",X"60",X"11",X"35",
		X"06",X"28",X"02",X"1E",X"B5",X"FF",X"3A",X"EF",X"89",X"A7",X"C8",X"CD",X"12",X"79",X"21",X"D1",
		X"15",X"E5",X"3A",X"0A",X"88",X"E6",X"1F",X"EF",X"01",X"16",X"B7",X"16",X"5D",X"17",X"C1",X"17",
		X"AF",X"18",X"EE",X"19",X"01",X"1A",X"64",X"1A",X"43",X"1B",X"8C",X"1B",X"AB",X"1B",X"CC",X"1B",
		X"03",X"1C",X"53",X"1C",X"66",X"1C",X"9C",X"1D",X"6E",X"1D",X"B2",X"6B",X"B9",X"71",X"FF",X"FF",
		X"FF",X"3A",X"06",X"88",X"A7",X"C0",X"3A",X"2C",X"88",X"FE",X"0F",X"CA",X"B5",X"0B",X"3A",X"02",
		X"88",X"A7",X"C8",X"21",X"05",X"88",X"36",X"02",X"2E",X"0A",X"36",X"00",X"CD",X"27",X"25",X"CD",
		X"B9",X"02",X"21",X"5F",X"85",X"11",X"E0",X"FF",X"06",X"08",X"3E",X"10",X"77",X"19",X"10",X"FA",
		X"C9",X"CD",X"C9",X"02",X"C0",X"CD",X"E3",X"02",X"CD",X"BC",X"19",X"AF",X"32",X"21",X"8D",X"21",
		X"23",X"8D",X"06",X"C0",X"D7",X"21",X"21",X"8E",X"06",X"0C",X"D7",X"32",X"16",X"8F",X"32",X"17",
		X"8F",X"3A",X"0E",X"88",X"A7",X"3E",X"02",X"28",X"2A",X"3A",X"E3",X"89",X"A7",X"20",X"24",X"3C",
		X"32",X"E3",X"89",X"3A",X"0F",X"88",X"A7",X"3A",X"0D",X"88",X"20",X"06",X"3D",X"32",X"1F",X"88",
		X"18",X"01",X"3D",X"11",X"02",X"06",X"A7",X"20",X"01",X"1C",X"FF",X"01",X"79",X"07",X"CD",X"5D",
		X"07",X"3E",X"80",X"32",X"08",X"88",X"21",X"0A",X"88",X"34",X"3A",X"0D",X"88",X"21",X"40",X"89",
		X"11",X"00",X"89",X"01",X"3F",X"00",X"A7",X"28",X"03",X"21",X"80",X"89",X"ED",X"B0",X"3A",X"03",
		X"89",X"A7",X"28",X"05",X"D6",X"02",X"32",X"31",X"89",X"3A",X"06",X"89",X"A7",X"C0",X"32",X"05",
		X"89",X"32",X"0A",X"89",X"11",X"AE",X"16",X"21",X"F0",X"89",X"1A",X"FE",X"FF",X"C8",X"77",X"13",
		X"23",X"18",X"F7",X"C9",X"11",X"AE",X"16",X"21",X"F0",X"89",X"1A",X"FE",X"FF",X"28",X"07",X"BE",
		X"20",X"15",X"13",X"23",X"18",X"F4",X"21",X"F0",X"89",X"AF",X"06",X"07",X"D7",X"C9",X"0A",X"10",
		X"1B",X"1F",X"1E",X"11",X"1D",X"19",X"FF",X"21",X"08",X"88",X"35",X"C0",X"CD",X"E3",X"02",X"CD",
		X"D3",X"1D",X"3A",X"50",X"8F",X"E6",X"01",X"28",X"06",X"3E",X"10",X"32",X"0A",X"88",X"C9",X"AF",
		X"32",X"B7",X"88",X"CD",X"C2",X"03",X"3A",X"50",X"8F",X"A7",X"28",X"17",X"3A",X"07",X"89",X"CB",
		X"4F",X"20",X"08",X"21",X"81",X"4E",X"11",X"39",X"50",X"18",X"3D",X"21",X"92",X"4C",X"11",X"CE",
		X"4D",X"18",X"35",X"3A",X"04",X"89",X"A7",X"20",X"1C",X"3A",X"06",X"88",X"A7",X"28",X"16",X"3A",
		X"07",X"89",X"CB",X"47",X"21",X"2C",X"46",X"11",X"30",X"4B",X"20",X"1C",X"A7",X"21",X"A9",X"44",
		X"11",X"55",X"4B",X"28",X"13",X"3A",X"07",X"89",X"CB",X"47",X"21",X"D6",X"46",X"11",X"50",X"4A",
		X"28",X"06",X"21",X"72",X"48",X"11",X"F6",X"4B",X"ED",X"53",X"45",X"8F",X"22",X"BA",X"88",X"21",
		X"42",X"84",X"22",X"B8",X"88",X"21",X"42",X"80",X"22",X"43",X"8F",X"3E",X"20",X"32",X"07",X"8D",
		X"21",X"0A",X"88",X"34",X"11",X"83",X"06",X"FF",X"CD",X"94",X"16",X"C9",X"FF",X"FF",X"E0",X"B0",
		X"80",X"40",X"20",X"00",X"04",X"08",X"8D",X"8F",X"0F",X"88",X"8E",X"8C",X"5A",X"CD",X"81",X"43",
		X"21",X"B7",X"88",X"34",X"7E",X"FE",X"1C",X"C0",X"36",X"00",X"21",X"20",X"89",X"7E",X"34",X"A7",
		X"C8",X"AF",X"77",X"3A",X"50",X"8F",X"A7",X"20",X"42",X"3A",X"04",X"89",X"A7",X"20",X"22",X"3A",
		X"06",X"88",X"A7",X"28",X"13",X"3A",X"07",X"89",X"CB",X"47",X"20",X"06",X"3A",X"07",X"89",X"A7",
		X"20",X"06",X"3E",X"0D",X"32",X"0A",X"88",X"C9",X"3E",X"01",X"32",X"04",X"89",X"3C",X"32",X"03",
		X"89",X"CD",X"AD",X"1E",X"CD",X"65",X"20",X"CD",X"0B",X"4A",X"3E",X"10",X"32",X"91",X"8A",X"32",
		X"06",X"8F",X"32",X"09",X"8F",X"CD",X"0D",X"54",X"CD",X"EF",X"02",X"21",X"0A",X"88",X"36",X"03",
		X"C9",X"DD",X"21",X"80",X"8A",X"3A",X"50",X"8F",X"A7",X"11",X"F6",X"84",X"20",X"0A",X"3A",X"07",
		X"89",X"CB",X"47",X"21",X"2C",X"1E",X"20",X"05",X"21",X"34",X"1E",X"1E",X"E9",X"ED",X"53",X"BE",
		X"88",X"11",X"18",X"00",X"06",X"04",X"DD",X"36",X"00",X"01",X"7E",X"DD",X"77",X"04",X"23",X"7E",
		X"DD",X"77",X"06",X"23",X"DD",X"19",X"10",X"EE",X"DD",X"21",X"80",X"8A",X"3A",X"1F",X"88",X"A7",
		X"20",X"06",X"DD",X"35",X"06",X"DD",X"35",X"06",X"21",X"C9",X"26",X"22",X"00",X"8F",X"CD",X"B1",
		X"22",X"3A",X"50",X"8F",X"A7",X"20",X"31",X"3A",X"06",X"88",X"A7",X"20",X"0C",X"3A",X"3F",X"8F",
		X"A7",X"28",X"06",X"21",X"0A",X"88",X"36",X"12",X"C9",X"21",X"0A",X"88",X"34",X"11",X"3F",X"18",
		X"21",X"F0",X"89",X"1A",X"FE",X"43",X"C8",X"D6",X"88",X"77",X"13",X"23",X"18",X"F5",X"C9",X"92",
		X"98",X"A3",X"A7",X"A6",X"99",X"A5",X"A1",X"43",X"3A",X"07",X"89",X"CB",X"4F",X"28",X"5A",X"3A",
		X"07",X"89",X"CB",X"3F",X"FE",X"07",X"38",X"06",X"3E",X"08",X"06",X"03",X"18",X"07",X"CB",X"3F",
		X"E6",X"03",X"47",X"C6",X"05",X"32",X"47",X"8F",X"78",X"21",X"EB",X"70",X"CD",X"45",X"0C",X"EB",
		X"DD",X"21",X"E0",X"8A",X"3A",X"47",X"8F",X"47",X"0E",X"00",X"DD",X"36",X"05",X"80",X"DD",X"36",
		X"00",X"01",X"DD",X"36",X"06",X"04",X"DD",X"74",X"04",X"7D",X"E6",X"0F",X"84",X"67",X"7D",X"E6",
		X"F0",X"81",X"4F",X"DD",X"77",X"03",X"30",X"04",X"DD",X"34",X"04",X"24",X"11",X"29",X"38",X"CD",
		X"1E",X"38",X"11",X"18",X"00",X"DD",X"19",X"10",X"D1",X"21",X"0A",X"88",X"36",X"0F",X"C9",X"CD",
		X"55",X"1E",X"CD",X"AB",X"6C",X"CD",X"D4",X"20",X"CD",X"1B",X"51",X"CD",X"77",X"33",X"CD",X"BD",
		X"40",X"CD",X"EF",X"02",X"CD",X"DA",X"18",X"CD",X"1C",X"19",X"CD",X"E4",X"5A",X"CD",X"6E",X"19",
		X"CD",X"2F",X"1F",X"CD",X"3B",X"6B",X"CD",X"CA",X"19",X"C9",X"3A",X"09",X"89",X"A7",X"28",X"2E",
		X"4F",X"3A",X"0D",X"88",X"21",X"A4",X"88",X"A7",X"28",X"03",X"21",X"A7",X"88",X"7E",X"B9",X"C0",
		X"21",X"08",X"89",X"7E",X"FE",X"FF",X"30",X"01",X"34",X"3A",X"00",X"88",X"A7",X"3E",X"08",X"28",
		X"01",X"3D",X"81",X"27",X"32",X"09",X"89",X"CD",X"C2",X"03",X"CD",X"0D",X"0F",X"C9",X"3A",X"00",
		X"88",X"A7",X"3E",X"05",X"28",X"02",X"3E",X"03",X"32",X"09",X"89",X"C9",X"3A",X"01",X"89",X"A7",
		X"C0",X"3A",X"82",X"8A",X"A7",X"C0",X"21",X"E2",X"8A",X"11",X"18",X"00",X"06",X"06",X"3E",X"03",
		X"BE",X"C8",X"19",X"10",X"FB",X"21",X"0A",X"88",X"34",X"3A",X"07",X"89",X"CB",X"47",X"20",X"15",
		X"CB",X"3F",X"47",X"3A",X"20",X"88",X"80",X"47",X"3A",X"03",X"89",X"80",X"47",X"FE",X"20",X"38",
		X"02",X"3E",X"1F",X"18",X"0B",X"47",X"3A",X"20",X"88",X"80",X"FE",X"20",X"38",X"02",X"3E",X"1F",
		X"32",X"00",X"89",X"AF",X"32",X"87",X"8A",X"32",X"05",X"89",X"32",X"06",X"89",X"C9",X"3A",X"55",
		X"8D",X"A7",X"C0",X"3A",X"02",X"89",X"FE",X"05",X"38",X"26",X"28",X"0E",X"32",X"55",X"8D",X"3A",
		X"32",X"8D",X"A7",X"20",X"03",X"CD",X"6C",X"0F",X"18",X"16",X"3A",X"32",X"8D",X"A7",X"20",X"03",
		X"21",X"68",X"8D",X"7E",X"A7",X"20",X"09",X"36",X"01",X"2C",X"2C",X"36",X"01",X"CD",X"58",X"0F",
		X"3A",X"21",X"8D",X"A7",X"C0",X"3A",X"24",X"8F",X"A7",X"C0",X"21",X"22",X"8D",X"7E",X"A7",X"28",
		X"02",X"35",X"C9",X"36",X"20",X"2D",X"36",X"01",X"CD",X"76",X"0F",X"C9",X"21",X"80",X"8A",X"11",
		X"81",X"8A",X"01",X"FF",X"01",X"36",X"00",X"ED",X"B0",X"C9",X"3A",X"06",X"88",X"A7",X"C0",X"3A",
		X"68",X"8D",X"A7",X"C8",X"21",X"6A",X"8D",X"35",X"C0",X"36",X"18",X"2D",X"CB",X"46",X"20",X"07",
		X"36",X"01",X"11",X"0F",X"06",X"FF",X"C9",X"36",X"00",X"11",X"8F",X"06",X"FF",X"C9",X"CD",X"8B",
		X"30",X"CD",X"A6",X"25",X"CD",X"77",X"33",X"CD",X"BD",X"40",X"CD",X"C6",X"28",X"CD",X"EF",X"02",
		X"C9",X"CD",X"27",X"25",X"32",X"02",X"89",X"32",X"34",X"89",X"0E",X"30",X"3A",X"07",X"89",X"FE",
		X"02",X"30",X"02",X"0E",X"28",X"21",X"01",X"89",X"71",X"2E",X"07",X"34",X"7E",X"E6",X"01",X"20",
		X"26",X"3A",X"06",X"88",X"A7",X"CA",X"3C",X"1D",X"3A",X"50",X"8F",X"A7",X"20",X"10",X"35",X"3E",
		X"01",X"32",X"50",X"8F",X"32",X"01",X"89",X"3E",X"40",X"32",X"4A",X"8F",X"18",X"09",X"AF",X"21",
		X"45",X"8F",X"06",X"10",X"D7",X"26",X"81",X"2E",X"04",X"36",X"00",X"11",X"40",X"89",X"21",X"00",
		X"89",X"01",X"3F",X"00",X"3A",X"0D",X"88",X"A7",X"28",X"03",X"11",X"80",X"89",X"ED",X"B0",X"AF",
		X"32",X"0A",X"88",X"C9",X"3A",X"50",X"8F",X"A7",X"20",X"97",X"CD",X"4E",X"0F",X"CD",X"27",X"25",
		X"AF",X"32",X"E3",X"89",X"3A",X"06",X"88",X"A7",X"CA",X"3C",X"1D",X"21",X"08",X"89",X"7E",X"A7",
		X"28",X"14",X"35",X"28",X"11",X"CD",X"C2",X"03",X"0E",X"0A",X"3A",X"0D",X"88",X"A7",X"28",X"01",
		X"0C",X"79",X"32",X"0A",X"88",X"C9",X"CD",X"92",X"0F",X"21",X"0A",X"88",X"3A",X"0D",X"88",X"A7",
		X"28",X"01",X"34",X"34",X"AF",X"32",X"FC",X"89",X"32",X"31",X"89",X"32",X"32",X"89",X"CD",X"B2",
		X"1A",X"C9",X"01",X"1E",X"00",X"68",X"11",X"03",X"00",X"DD",X"21",X"A2",X"88",X"3A",X"0D",X"88",
		X"0F",X"30",X"02",X"DD",X"19",X"FD",X"21",X"00",X"8A",X"DD",X"7E",X"02",X"FD",X"BE",X"02",X"20",
		X"0E",X"DD",X"7E",X"01",X"FD",X"BE",X"01",X"20",X"06",X"DD",X"7E",X"00",X"FD",X"BE",X"00",X"30",
		X"09",X"FD",X"19",X"2C",X"0D",X"0D",X"0D",X"C8",X"18",X"DF",X"7D",X"3C",X"32",X"FC",X"89",X"3D",
		X"C5",X"21",X"1D",X"8A",X"11",X"20",X"8A",X"ED",X"B8",X"6F",X"DD",X"7E",X"00",X"FD",X"77",X"00",
		X"DD",X"7E",X"01",X"FD",X"77",X"01",X"DD",X"7E",X"02",X"FD",X"77",X"02",X"C1",X"C5",X"DD",X"21",
		X"30",X"8A",X"21",X"E1",X"89",X"3A",X"0D",X"88",X"A7",X"28",X"05",X"DD",X"21",X"33",X"8A",X"23",
		X"36",X"01",X"2E",X"DD",X"11",X"E0",X"89",X"ED",X"B8",X"DD",X"7E",X"02",X"12",X"1B",X"DD",X"7E",
		X"01",X"12",X"C1",X"21",X"1C",X"8E",X"11",X"1F",X"8E",X"ED",X"B8",X"EB",X"2B",X"3E",X"10",X"06",
		X"03",X"D7",X"C9",X"CD",X"C9",X"02",X"C0",X"CD",X"E3",X"02",X"01",X"19",X"08",X"CD",X"5D",X"07",
		X"11",X"00",X"06",X"FF",X"1E",X"02",X"FF",X"CD",X"60",X"79",X"3E",X"0C",X"32",X"0A",X"88",X"AF",
		X"32",X"08",X"88",X"11",X"93",X"55",X"01",X"00",X"22",X"1A",X"E6",X"37",X"0F",X"89",X"4F",X"13",
		X"10",X"F7",X"FE",X"7C",X"28",X"04",X"21",X"1E",X"88",X"34",X"11",X"F2",X"1F",X"21",X"F0",X"89",
		X"1A",X"FE",X"A0",X"C8",X"C6",X"08",X"77",X"13",X"23",X"18",X"F5",X"C9",X"CD",X"C9",X"02",X"C0",
		X"01",X"19",X"08",X"CD",X"5D",X"07",X"11",X"00",X"06",X"FF",X"1E",X"03",X"FF",X"CD",X"60",X"79",
		X"3E",X"0C",X"32",X"0A",X"88",X"3E",X"60",X"32",X"08",X"88",X"C9",X"3A",X"0E",X"88",X"A7",X"28",
		X"0B",X"3A",X"88",X"89",X"A7",X"28",X"05",X"3E",X"01",X"32",X"0D",X"88",X"11",X"40",X"89",X"21",
		X"00",X"89",X"01",X"3F",X"00",X"ED",X"B0",X"AF",X"32",X"0A",X"88",X"C9",X"3A",X"48",X"89",X"A7",
		X"28",X"04",X"AF",X"32",X"0D",X"88",X"11",X"80",X"89",X"21",X"00",X"89",X"01",X"3F",X"00",X"ED",
		X"B0",X"AF",X"32",X"0A",X"88",X"21",X"28",X"53",X"06",X"0E",X"7E",X"E6",X"1F",X"83",X"5F",X"30",
		X"01",X"14",X"23",X"10",X"F5",X"3E",X"60",X"BB",X"20",X"04",X"3E",X"8A",X"92",X"C8",X"21",X"38",
		X"8A",X"34",X"C9",X"21",X"08",X"88",X"35",X"C0",X"3E",X"82",X"CD",X"B2",X"05",X"3E",X"80",X"CD",
		X"B2",X"05",X"3E",X"89",X"CD",X"B2",X"05",X"01",X"D9",X"07",X"CD",X"5D",X"07",X"CD",X"E9",X"03",
		X"11",X"11",X"06",X"FF",X"21",X"0A",X"88",X"36",X"0E",X"3A",X"FC",X"89",X"A7",X"C8",X"21",X"45",
		X"80",X"47",X"2C",X"2C",X"10",X"FC",X"22",X"FD",X"89",X"CD",X"C1",X"0F",X"21",X"FF",X"89",X"36",
		X"07",X"11",X"54",X"17",X"21",X"F0",X"89",X"1A",X"FE",X"5A",X"C8",X"CB",X"17",X"77",X"13",X"23",
		X"18",X"F5",X"C9",X"3A",X"07",X"89",X"E6",X"01",X"20",X"05",X"CD",X"E2",X"64",X"18",X"03",X"CD",
		X"F8",X"68",X"CD",X"EF",X"02",X"C9",X"21",X"08",X"88",X"35",X"3A",X"2A",X"8E",X"A7",X"28",X"04",
		X"7E",X"A7",X"28",X"28",X"CD",X"94",X"7E",X"3A",X"FC",X"89",X"A7",X"C8",X"3A",X"08",X"88",X"E6",
		X"07",X"C0",X"3A",X"FF",X"89",X"2A",X"FD",X"89",X"11",X"20",X"00",X"06",X"1C",X"77",X"19",X"10",
		X"FC",X"3C",X"FE",X"10",X"38",X"02",X"3E",X"06",X"32",X"FF",X"89",X"C9",X"21",X"5F",X"85",X"11",
		X"E0",X"FF",X"06",X"08",X"3E",X"10",X"77",X"19",X"10",X"FA",X"21",X"BC",X"82",X"11",X"E0",X"FF",
		X"01",X"00",X"0A",X"7E",X"81",X"4F",X"19",X"10",X"FA",X"79",X"FE",X"AA",X"C0",X"AF",X"32",X"2A",
		X"8E",X"3A",X"0E",X"88",X"A7",X"28",X"4E",X"3A",X"0D",X"88",X"A7",X"28",X"29",X"3A",X"48",X"89",
		X"A7",X"28",X"42",X"AF",X"32",X"0D",X"88",X"32",X"0A",X"88",X"21",X"80",X"89",X"06",X"3F",X"D7",
		X"3C",X"32",X"1F",X"88",X"CD",X"E3",X"02",X"21",X"E0",X"84",X"36",X"02",X"11",X"E0",X"FF",X"19",
		X"36",X"25",X"19",X"36",X"20",X"C9",X"3A",X"88",X"89",X"A7",X"28",X"19",X"AF",X"32",X"0A",X"88",
		X"21",X"40",X"89",X"06",X"3F",X"D7",X"3C",X"32",X"0D",X"88",X"CD",X"E3",X"02",X"21",X"40",X"87",
		X"36",X"01",X"18",X"D8",X"C9",X"AF",X"21",X"00",X"89",X"06",X"BF",X"D7",X"3A",X"0E",X"88",X"A7",
		X"CC",X"0D",X"1D",X"C4",X"E7",X"1C",X"3A",X"02",X"88",X"A7",X"28",X"10",X"AF",X"32",X"06",X"88",
		X"32",X"0A",X"88",X"3C",X"32",X"1F",X"88",X"3C",X"32",X"05",X"88",X"C9",X"AF",X"32",X"06",X"88",
		X"32",X"0A",X"88",X"32",X"0D",X"88",X"32",X"0E",X"88",X"32",X"51",X"8E",X"3C",X"32",X"05",X"88",
		X"32",X"1F",X"88",X"32",X"3F",X"8F",X"CD",X"B9",X"02",X"CD",X"CF",X"0E",X"11",X"4C",X"1E",X"21",
		X"F0",X"89",X"1A",X"FE",X"7F",X"C8",X"CB",X"3F",X"77",X"13",X"23",X"18",X"F5",X"C9",X"21",X"4A",
		X"8F",X"7E",X"35",X"FE",X"40",X"20",X"0B",X"CD",X"E9",X"79",X"11",X"26",X"06",X"FF",X"CD",X"44",
		X"0F",X"C9",X"A7",X"C0",X"32",X"0A",X"88",X"2E",X"50",X"36",X"02",X"21",X"07",X"8D",X"36",X"40",
		X"3A",X"07",X"89",X"CB",X"4F",X"C0",X"3E",X"01",X"32",X"61",X"8F",X"C9",X"3A",X"07",X"89",X"CB",
		X"4F",X"20",X"04",X"CD",X"D5",X"0F",X"C9",X"CD",X"A6",X"6D",X"21",X"4C",X"58",X"7D",X"D6",X"24",
		X"6F",X"24",X"24",X"01",X"20",X"20",X"AF",X"CB",X"46",X"28",X"01",X"3C",X"CB",X"5E",X"20",X"01",
		X"3C",X"10",X"F4",X"B9",X"C8",X"3E",X"01",X"32",X"E7",X"89",X"C9",X"10",X"12",X"14",X"18",X"1A",
		X"1C",X"1E",X"20",X"3A",X"04",X"89",X"A7",X"21",X"07",X"89",X"20",X"0F",X"3A",X"06",X"88",X"A7",
		X"28",X"09",X"7E",X"CB",X"47",X"20",X"2A",X"7E",X"A7",X"28",X"26",X"7E",X"E6",X"01",X"01",X"39",
		X"08",X"20",X"03",X"01",X"79",X"08",X"CD",X"5D",X"07",X"3E",X"0F",X"21",X"45",X"80",X"11",X"20",
		X"00",X"06",X"04",X"77",X"19",X"10",X"FC",X"21",X"46",X"80",X"06",X"04",X"77",X"19",X"10",X"FC",
		X"C9",X"3A",X"50",X"8F",X"A7",X"20",X"D4",X"01",X"59",X"08",X"CD",X"5D",X"07",X"21",X"1C",X"81",
		X"11",X"20",X"00",X"06",X"10",X"3E",X"09",X"77",X"19",X"10",X"FC",X"C9",X"C0",X"B0",X"BA",X"00",
		X"B0",X"C0",X"C0",X"C0",X"58",X"B0",X"52",X"00",X"48",X"C0",X"58",X"C0",X"05",X"04",X"03",X"03",
		X"02",X"01",X"01",X"00",X"08",X"07",X"06",X"05",X"04",X"03",X"02",X"01",X"14",X"30",X"36",X"3E",
		X"3C",X"22",X"3A",X"32",X"7F",X"21",X"E5",X"89",X"46",X"7D",X"C6",X"16",X"6F",X"78",X"B6",X"A7",
		X"DD",X"21",X"80",X"8A",X"20",X"3C",X"3A",X"06",X"88",X"A7",X"C8",X"FD",X"21",X"90",X"8C",X"DD",
		X"7E",X"02",X"A7",X"20",X"2D",X"3A",X"24",X"8F",X"21",X"57",X"8F",X"B6",X"20",X"24",X"3A",X"1F",
		X"88",X"A7",X"3A",X"A0",X"A0",X"20",X"03",X"3A",X"C0",X"A0",X"2F",X"DD",X"77",X"07",X"17",X"17",
		X"17",X"21",X"03",X"8F",X"17",X"CB",X"16",X"7E",X"E6",X"07",X"FE",X"01",X"C8",X"DD",X"CB",X"07",
		X"A6",X"C9",X"DD",X"36",X"07",X"00",X"C9",X"22",X"1F",X"25",X"1E",X"14",X"10",X"3A",X"1E",X"88",
		X"A7",X"20",X"5E",X"21",X"5F",X"85",X"01",X"A7",X"1E",X"11",X"E0",X"FF",X"0A",X"77",X"03",X"19",
		X"FE",X"10",X"20",X"F8",X"3A",X"07",X"89",X"3C",X"47",X"AF",X"C6",X"01",X"27",X"10",X"FB",X"F5",
		X"F5",X"F5",X"CB",X"3F",X"CB",X"3F",X"CB",X"3F",X"CB",X"3F",X"21",X"9F",X"84",X"A7",X"20",X"02",
		X"3E",X"10",X"77",X"F1",X"E6",X"0F",X"21",X"7F",X"84",X"77",X"F1",X"CB",X"3F",X"CB",X"3F",X"CB",
		X"3F",X"CB",X"3F",X"E6",X"01",X"21",X"0D",X"20",X"CD",X"45",X"0C",X"21",X"62",X"84",X"CD",X"07",
		X"33",X"21",X"22",X"87",X"CD",X"8C",X"1F",X"F1",X"47",X"E6",X"0F",X"32",X"83",X"84",X"CD",X"FB",
		X"1F",X"CD",X"18",X"1F",X"CD",X"C9",X"34",X"C9",X"21",X"E7",X"89",X"06",X"07",X"7E",X"23",X"B6",
		X"C0",X"10",X"FA",X"0E",X"00",X"2E",X"01",X"7E",X"D6",X"0A",X"38",X"22",X"0C",X"18",X"F9",X"3A",
		X"56",X"8D",X"A7",X"C0",X"4F",X"3A",X"01",X"89",X"FE",X"0A",X"38",X"0D",X"21",X"87",X"1F",X"06",
		X"05",X"BE",X"28",X"0A",X"0C",X"23",X"10",X"F9",X"C9",X"3E",X"01",X"32",X"56",X"8D",X"79",X"A7",
		X"20",X"28",X"3A",X"07",X"89",X"C6",X"01",X"47",X"AF",X"C6",X"01",X"27",X"10",X"FB",X"11",X"E6",
		X"1F",X"CB",X"67",X"20",X"03",X"11",X"DA",X"1F",X"21",X"22",X"87",X"CD",X"8C",X"1F",X"3E",X"10",
		X"06",X"03",X"D7",X"3A",X"01",X"89",X"32",X"43",X"87",X"AF",X"21",X"A3",X"1F",X"CD",X"45",X"0C",
		X"21",X"22",X"83",X"CD",X"8C",X"1F",X"C9",X"09",X"14",X"1E",X"28",X"30",X"3E",X"04",X"ED",X"47",
		X"06",X"03",X"1A",X"77",X"2C",X"13",X"10",X"FA",X"0E",X"1D",X"09",X"ED",X"57",X"3D",X"C8",X"ED",
		X"47",X"18",X"ED",X"AD",X"1F",X"B6",X"1F",X"C2",X"1F",X"CE",X"1F",X"44",X"20",X"8E",X"8E",X"8E",
		X"8E",X"00",X"CE",X"8E",X"8E",X"CE",X"8F",X"8F",X"8F",X"8F",X"00",X"CF",X"8F",X"00",X"CF",X"0F",
		X"0F",X"0F",X"85",X"85",X"85",X"85",X"00",X"C5",X"85",X"00",X"C5",X"05",X"05",X"05",X"8B",X"8B",
		X"8B",X"8B",X"00",X"CB",X"8B",X"00",X"CB",X"0B",X"0B",X"0B",X"B7",X"B8",X"B9",X"B6",X"09",X"B6",
		X"B2",X"B3",X"B2",X"10",X"10",X"10",X"B7",X"B8",X"B9",X"B6",X"09",X"B6",X"B4",X"B5",X"B4",X"10",
		X"10",X"10",X"02",X"08",X"13",X"17",X"16",X"09",X"15",X"11",X"A0",X"78",X"CB",X"6F",X"11",X"3B",
		X"20",X"28",X"03",X"11",X"50",X"20",X"21",X"62",X"80",X"CD",X"07",X"33",X"C9",X"11",X"20",X"26",
		X"20",X"B2",X"B3",X"B2",X"B6",X"10",X"B6",X"B7",X"B8",X"B9",X"B7",X"B8",X"B9",X"B6",X"B1",X"B6",
		X"B6",X"10",X"B6",X"B7",X"B8",X"B9",X"B4",X"B5",X"B4",X"B6",X"10",X"B6",X"B7",X"B8",X"B9",X"B7",
		X"B8",X"B9",X"B6",X"B1",X"B6",X"B6",X"10",X"B6",X"B7",X"B8",X"B9",X"00",X"00",X"40",X"00",X"00",
		X"40",X"00",X"00",X"00",X"83",X"83",X"83",X"83",X"00",X"C3",X"83",X"00",X"C3",X"03",X"03",X"03",
		X"0B",X"0B",X"4B",X"0B",X"00",X"4B",X"0B",X"0B",X"0B",X"83",X"83",X"83",X"83",X"00",X"C3",X"83",
		X"00",X"C3",X"03",X"03",X"03",X"21",X"3F",X"86",X"11",X"E0",X"FF",X"3A",X"08",X"89",X"A7",X"C8",
		X"3D",X"4F",X"28",X"0D",X"FE",X"05",X"38",X"02",X"3E",X"05",X"4F",X"47",X"36",X"B0",X"19",X"10",
		X"FB",X"3E",X"05",X"91",X"C8",X"47",X"36",X"10",X"19",X"10",X"FB",X"C9",X"21",X"6D",X"06",X"06",
		X"10",X"11",X"AA",X"20",X"1A",X"BE",X"20",X"0C",X"13",X"00",X"3E",X"08",X"85",X"30",X"01",X"24",
		X"6F",X"10",X"F1",X"C9",X"3E",X"01",X"32",X"F0",X"8E",X"C9",X"F5",X"D5",X"80",X"94",X"88",X"18",
		X"03",X"0B",X"06",X"15",X"32",X"88",X"77",X"3A",X"35",X"CD",X"05",X"0C",X"32",X"D1",X"3E",X"DD",
		X"2C",X"2C",X"0A",X"10",X"1B",X"1F",X"1E",X"11",X"1D",X"19",X"FF",X"00",X"00",X"00",X"11",X"00",
		X"0E",X"00",X"00",X"07",X"21",X"32",X"8D",X"3A",X"50",X"8F",X"A7",X"28",X"0B",X"36",X"00",X"45",
		X"2E",X"F8",X"7E",X"23",X"A6",X"20",X"03",X"68",X"7E",X"A7",X"C2",X"1E",X"24",X"DD",X"21",X"80",
		X"8A",X"CD",X"29",X"23",X"CD",X"01",X"21",X"CD",X"63",X"25",X"CD",X"A6",X"25",X"CD",X"8B",X"30",
		X"C9",X"CD",X"78",X"27",X"CD",X"0B",X"21",X"CD",X"57",X"21",X"C9",X"DD",X"21",X"80",X"8A",X"DD",
		X"CB",X"07",X"66",X"DD",X"36",X"07",X"00",X"C8",X"21",X"02",X"8F",X"7E",X"A7",X"C0",X"34",X"FD",
		X"21",X"90",X"8C",X"3A",X"30",X"8F",X"FE",X"02",X"38",X"15",X"FD",X"7E",X"18",X"FE",X"02",X"20",
		X"0E",X"FD",X"7E",X"00",X"A7",X"20",X"08",X"FD",X"36",X"18",X"00",X"FD",X"CB",X"00",X"CE",X"11",
		X"18",X"00",X"06",X"02",X"FD",X"CB",X"00",X"46",X"28",X"3A",X"FD",X"19",X"10",X"F6",X"DD",X"54",
		X"1E",X"3C",X"1A",X"A7",X"20",X"01",X"C9",X"FD",X"21",X"90",X"8C",X"3E",X"02",X"32",X"15",X"8F",
		X"FD",X"CB",X"00",X"46",X"C4",X"CF",X"21",X"11",X"18",X"00",X"FD",X"19",X"3A",X"15",X"8F",X"D6",
		X"01",X"20",X"EA",X"3A",X"00",X"8F",X"11",X"C9",X"26",X"D6",X"0C",X"93",X"C2",X"B1",X"22",X"AF",
		X"32",X"02",X"8F",X"C9",X"FD",X"CB",X"00",X"C6",X"DD",X"7E",X"04",X"D6",X"03",X"FD",X"77",X"04",
		X"DD",X"7E",X"06",X"C6",X"04",X"FD",X"77",X"06",X"FD",X"CB",X"00",X"4E",X"20",X"0A",X"FD",X"36",
		X"0F",X"14",X"FD",X"36",X"10",X"40",X"18",X"14",X"FD",X"36",X"0F",X"10",X"FD",X"36",X"10",X"40",
		X"3E",X"01",X"32",X"77",X"8D",X"AF",X"21",X"98",X"8A",X"06",X"18",X"D7",X"21",X"19",X"8D",X"FD",
		X"E5",X"D1",X"AF",X"CB",X"5B",X"28",X"01",X"23",X"77",X"23",X"23",X"77",X"C3",X"B1",X"22",X"FD",
		X"CB",X"07",X"46",X"20",X"2F",X"FD",X"7E",X"12",X"A7",X"20",X"06",X"FD",X"34",X"12",X"CD",X"D2",
		X"0E",X"FD",X"CB",X"00",X"4E",X"20",X"3F",X"FD",X"7D",X"CB",X"5F",X"21",X"1B",X"8D",X"28",X"01",
		X"23",X"7E",X"A7",X"28",X"04",X"36",X"00",X"18",X"25",X"FD",X"7E",X"06",X"D6",X"04",X"38",X"1E",
		X"FD",X"77",X"06",X"C9",X"FD",X"7E",X"01",X"FE",X"01",X"D8",X"20",X"07",X"FD",X"36",X"0F",X"1B",
		X"FD",X"34",X"01",X"FD",X"7E",X"04",X"C6",X"04",X"FD",X"77",X"04",X"FE",X"E8",X"D8",X"FD",X"E5",
		X"E1",X"06",X"18",X"AF",X"D7",X"C9",X"3A",X"0E",X"8F",X"A7",X"CC",X"82",X"22",X"ED",X"5B",X"10",
		X"8F",X"FD",X"7D",X"CB",X"5F",X"FD",X"6E",X"05",X"FD",X"66",X"06",X"01",X"19",X"8D",X"28",X"01",
		X"03",X"0A",X"CB",X"47",X"28",X"03",X"19",X"18",X"02",X"ED",X"52",X"FD",X"75",X"05",X"FD",X"74",
		X"06",X"ED",X"5B",X"12",X"8F",X"FD",X"6E",X"03",X"FD",X"66",X"04",X"19",X"7C",X"FE",X"E8",X"30",
		X"0B",X"FD",X"75",X"03",X"FD",X"74",X"04",X"21",X"0E",X"8F",X"35",X"C9",X"AF",X"32",X"0E",X"8F",
		X"32",X"0F",X"8F",X"32",X"30",X"8F",X"32",X"45",X"8D",X"32",X"77",X"8D",X"32",X"3F",X"8F",X"18",
		X"9D",X"C9",X"3A",X"0F",X"8F",X"21",X"12",X"27",X"E7",X"32",X"0E",X"8F",X"3A",X"0F",X"8F",X"21",
		X"1C",X"27",X"CD",X"45",X"0C",X"ED",X"53",X"10",X"8F",X"3A",X"0F",X"8F",X"21",X"30",X"27",X"CD",
		X"45",X"0C",X"ED",X"53",X"12",X"8F",X"21",X"0F",X"8F",X"34",X"7E",X"FE",X"09",X"C0",X"36",X"08",
		X"C9",X"3A",X"32",X"8D",X"A7",X"C0",X"DD",X"21",X"80",X"8A",X"CD",X"E6",X"22",X"11",X"18",X"00",
		X"DD",X"19",X"CD",X"E6",X"22",X"DD",X"19",X"CD",X"E6",X"22",X"DD",X"19",X"CD",X"E6",X"22",X"C9",
		X"FD",X"21",X"90",X"8C",X"11",X"18",X"00",X"06",X"02",X"AF",X"FD",X"CB",X"00",X"46",X"28",X"01",
		X"07",X"FD",X"19",X"10",X"F5",X"C9",X"DD",X"7E",X"0E",X"A7",X"28",X"04",X"DD",X"35",X"0E",X"C9",
		X"2A",X"00",X"8F",X"7E",X"FE",X"FF",X"28",X"12",X"DD",X"77",X"10",X"23",X"7E",X"DD",X"77",X"0F",
		X"23",X"7E",X"DD",X"77",X"0E",X"23",X"22",X"00",X"8F",X"C9",X"CD",X"D0",X"22",X"FE",X"03",X"20",
		X"08",X"21",X"E7",X"26",X"22",X"00",X"8F",X"18",X"D7",X"23",X"7E",X"32",X"00",X"8F",X"23",X"7E",
		X"32",X"01",X"8F",X"18",X"CB",X"10",X"10",X"37",X"37",X"DD",X"CB",X"07",X"56",X"28",X"3B",X"DD",
		X"35",X"04",X"DD",X"7E",X"04",X"FE",X"41",X"30",X"04",X"DD",X"36",X"04",X"41",X"CD",X"D7",X"23",
		X"2A",X"BE",X"88",X"7D",X"FE",X"E6",X"20",X"11",X"7E",X"FE",X"35",X"30",X"0C",X"26",X"89",X"06",
		X"07",X"23",X"7E",X"B7",X"20",X"03",X"10",X"F9",X"C9",X"CD",X"EC",X"23",X"21",X"BD",X"88",X"34",
		X"7E",X"E6",X"07",X"77",X"A7",X"C0",X"2B",X"34",X"18",X"43",X"DD",X"CB",X"07",X"5E",X"C8",X"DD",
		X"34",X"04",X"DD",X"7E",X"04",X"FE",X"C0",X"38",X"04",X"DD",X"36",X"04",X"C0",X"CD",X"D7",X"23",
		X"3A",X"BE",X"88",X"FE",X"F6",X"20",X"17",X"21",X"38",X"8A",X"06",X"03",X"7E",X"A7",X"20",X"0E",
		X"23",X"10",X"F9",X"21",X"83",X"80",X"3A",X"43",X"83",X"86",X"E6",X"0F",X"A7",X"C8",X"CD",X"05",
		X"24",X"21",X"BD",X"88",X"35",X"7E",X"E6",X"07",X"77",X"A7",X"C0",X"2B",X"35",X"7E",X"E6",X"03",
		X"77",X"21",X"F6",X"26",X"CD",X"45",X"0C",X"D5",X"21",X"25",X"84",X"CD",X"25",X"33",X"D1",X"2E",
		X"65",X"CD",X"25",X"33",X"2E",X"A5",X"11",X"0A",X"27",X"3A",X"BC",X"88",X"E6",X"01",X"20",X"03",
		X"11",X"0E",X"27",X"CD",X"25",X"33",X"C9",X"DD",X"21",X"80",X"8A",X"DD",X"7E",X"04",X"DD",X"77",
		X"4C",X"D6",X"10",X"DD",X"77",X"34",X"C6",X"0A",X"DD",X"77",X"1C",X"C9",X"21",X"37",X"8F",X"34",
		X"CB",X"46",X"C0",X"2A",X"BE",X"88",X"7E",X"FE",X"34",X"28",X"03",X"35",X"18",X"03",X"36",X"10",
		X"2B",X"22",X"BE",X"88",X"C9",X"21",X"37",X"8F",X"34",X"CB",X"46",X"C8",X"2A",X"BE",X"88",X"7E",
		X"FE",X"37",X"30",X"03",X"34",X"18",X"03",X"23",X"36",X"34",X"22",X"BE",X"88",X"C9",X"CD",X"01",
		X"21",X"CD",X"A6",X"25",X"CD",X"8B",X"30",X"3A",X"1E",X"88",X"A7",X"C0",X"DD",X"21",X"80",X"8A",
		X"DD",X"7E",X"02",X"E6",X"07",X"EF",X"42",X"24",X"73",X"24",X"97",X"24",X"B9",X"24",X"DB",X"24",
		X"FB",X"24",X"21",X"E8",X"89",X"7E",X"2E",X"EF",X"B6",X"C0",X"DD",X"36",X"11",X"10",X"DD",X"34",
		X"02",X"21",X"80",X"8A",X"11",X"98",X"8A",X"01",X"18",X"00",X"ED",X"B0",X"DD",X"7E",X"04",X"D6",
		X"10",X"DD",X"77",X"04",X"21",X"BD",X"26",X"CD",X"0F",X"25",X"3A",X"24",X"8F",X"A7",X"C0",X"CD",
		X"AD",X"0F",X"C9",X"DD",X"35",X"11",X"C0",X"3A",X"39",X"8A",X"A7",X"20",X"06",X"DD",X"36",X"11",
		X"10",X"DD",X"34",X"02",X"DD",X"7E",X"04",X"C6",X"10",X"DD",X"77",X"04",X"AF",X"DD",X"77",X"1E",
		X"21",X"C1",X"26",X"CD",X"0F",X"25",X"C9",X"DD",X"35",X"11",X"C0",X"DD",X"34",X"02",X"21",X"C5",
		X"26",X"CD",X"0F",X"25",X"DD",X"21",X"80",X"8A",X"DD",X"7E",X"04",X"C6",X"04",X"DD",X"77",X"04",
		X"DD",X"7E",X"06",X"D6",X"06",X"DD",X"77",X"06",X"C9",X"DD",X"34",X"05",X"DD",X"CB",X"05",X"46",
		X"20",X"03",X"DD",X"35",X"06",X"DD",X"7E",X"04",X"C6",X"02",X"DD",X"77",X"04",X"FE",X"DC",X"D8",
		X"CD",X"21",X"0F",X"DD",X"36",X"11",X"02",X"DD",X"34",X"02",X"C9",X"DD",X"35",X"11",X"C0",X"DD",
		X"7E",X"04",X"C6",X"04",X"DD",X"77",X"04",X"DD",X"7E",X"06",X"D6",X"08",X"DD",X"77",X"06",X"DD",
		X"36",X"0F",X"1A",X"DD",X"36",X"11",X"30",X"DD",X"34",X"02",X"C9",X"DD",X"35",X"11",X"C0",X"21",
		X"2B",X"88",X"7E",X"A7",X"20",X"02",X"2E",X"0A",X"36",X"07",X"3A",X"3C",X"8A",X"A7",X"C8",X"11",
		X"18",X"00",X"06",X"04",X"7E",X"DD",X"77",X"0F",X"23",X"DD",X"19",X"10",X"F7",X"21",X"E5",X"89",
		X"3A",X"F9",X"8D",X"B6",X"20",X"01",X"C9",X"16",X"08",X"FF",X"21",X"02",X"89",X"7E",X"FE",X"07",
		X"3E",X"00",X"38",X"0D",X"3A",X"FB",X"89",X"36",X"04",X"2E",X"34",X"36",X"04",X"06",X"20",X"68",
		X"D7",X"21",X"00",X"8F",X"06",X"4F",X"D7",X"2E",X"57",X"06",X"04",X"D7",X"21",X"30",X"8D",X"06",
		X"03",X"D7",X"32",X"82",X"8A",X"32",X"90",X"8C",X"32",X"A8",X"8C",X"32",X"52",X"8F",X"32",X"63",
		X"8F",X"C9",X"76",X"3A",X"50",X"8F",X"A7",X"C0",X"21",X"06",X"8F",X"7E",X"A7",X"28",X"02",X"35",
		X"C9",X"36",X"0C",X"23",X"34",X"EB",X"3A",X"07",X"89",X"CB",X"47",X"21",X"BB",X"87",X"1A",X"20",
		X"0E",X"26",X"84",X"11",X"44",X"27",X"E6",X"01",X"28",X"0F",X"11",X"48",X"27",X"18",X"0A",X"11",
		X"4C",X"27",X"E6",X"01",X"28",X"03",X"11",X"50",X"27",X"D5",X"CD",X"25",X"33",X"11",X"A0",X"FF",
		X"19",X"D1",X"CD",X"25",X"33",X"C9",X"3A",X"07",X"89",X"CB",X"47",X"CA",X"66",X"2D",X"21",X"09",
		X"8F",X"35",X"C0",X"36",X"10",X"3A",X"02",X"89",X"A7",X"C8",X"4F",X"3A",X"20",X"89",X"A7",X"20",
		X"74",X"79",X"11",X"05",X"8F",X"21",X"34",X"89",X"BE",X"28",X"10",X"1A",X"A7",X"20",X"0C",X"34",
		X"3C",X"12",X"11",X"E3",X"86",X"ED",X"53",X"32",X"89",X"18",X"10",X"1A",X"A7",X"28",X"0C",X"3A",
		X"32",X"89",X"FE",X"A3",X"20",X"05",X"AF",X"12",X"32",X"63",X"8F",X"7E",X"FE",X"07",X"38",X"0E",
		X"3A",X"32",X"89",X"FE",X"C3",X"20",X"05",X"3E",X"01",X"32",X"04",X"8F",X"3E",X"07",X"47",X"11",
		X"C0",X"FF",X"3A",X"05",X"8F",X"A7",X"28",X"63",X"21",X"09",X"8F",X"36",X"1C",X"11",X"E0",X"FF",
		X"DD",X"2A",X"32",X"89",X"DD",X"19",X"DD",X"22",X"32",X"89",X"23",X"CB",X"46",X"21",X"6C",X"27",
		X"20",X"03",X"21",X"68",X"27",X"DD",X"36",X"40",X"10",X"DD",X"36",X"41",X"10",X"CD",X"19",X"0F",
		X"CD",X"11",X"0F",X"18",X"43",X"3A",X"0A",X"8F",X"CB",X"47",X"21",X"70",X"27",X"28",X"03",X"21",
		X"74",X"27",X"FD",X"2A",X"32",X"89",X"FD",X"7C",X"D6",X"04",X"FD",X"67",X"FD",X"7E",X"00",X"FE",
		X"80",X"06",X"07",X"28",X"23",X"3E",X"80",X"11",X"C0",X"FF",X"FD",X"77",X"00",X"FD",X"77",X"01",
		X"FD",X"19",X"10",X"F6",X"CD",X"49",X"0F",X"06",X"07",X"18",X"0D",X"3A",X"0A",X"8F",X"CB",X"47",
		X"21",X"68",X"27",X"28",X"03",X"21",X"6C",X"27",X"DD",X"2A",X"32",X"89",X"11",X"C0",X"FF",X"E5",
		X"7E",X"DD",X"77",X"00",X"23",X"7E",X"DD",X"77",X"01",X"23",X"7E",X"DD",X"77",X"20",X"23",X"7E",
		X"DD",X"77",X"21",X"DD",X"19",X"E1",X"10",X"E7",X"3A",X"20",X"89",X"A7",X"20",X"1A",X"11",X"DF",
		X"FF",X"DD",X"19",X"DD",X"E5",X"E1",X"3A",X"0A",X"8F",X"CB",X"47",X"11",X"54",X"27",X"28",X"03",
		X"11",X"5E",X"27",X"CD",X"07",X"33",X"36",X"10",X"21",X"0A",X"8F",X"34",X"C9",X"05",X"08",X"0A",
		X"07",X"0C",X"10",X"0A",X"0F",X"0E",X"10",X"0A",X"0F",X"40",X"13",X"00",X"40",X"10",X"00",X"40",
		X"11",X"00",X"40",X"12",X"00",X"FF",X"D8",X"26",X"40",X"17",X"08",X"40",X"10",X"08",X"40",X"25",
		X"08",X"40",X"16",X"08",X"FF",X"E7",X"26",X"40",X"18",X"08",X"40",X"10",X"08",X"40",X"25",X"08",
		X"40",X"16",X"08",X"FF",X"C9",X"26",X"FE",X"26",X"02",X"27",X"FE",X"26",X"06",X"27",X"E8",X"E9",
		X"EB",X"EA",X"E4",X"E5",X"E7",X"E6",X"EC",X"ED",X"EF",X"EE",X"A8",X"A9",X"AB",X"AA",X"AC",X"AD",
		X"AB",X"AE",X"0B",X"04",X"08",X"08",X"0A",X"0A",X"08",X"08",X"08",X"18",X"00",X"03",X"C0",X"02",
		X"80",X"02",X"00",X"02",X"80",X"01",X"00",X"01",X"C0",X"00",X"80",X"00",X"40",X"00",X"00",X"00",
		X"00",X"00",X"40",X"00",X"80",X"00",X"C0",X"00",X"00",X"01",X"80",X"01",X"00",X"02",X"80",X"02",
		X"C0",X"02",X"00",X"03",X"3D",X"81",X"BD",X"42",X"5C",X"BF",X"BE",X"BB",X"D0",X"D1",X"D3",X"D2",
		X"D4",X"D5",X"D7",X"D6",X"10",X"C1",X"CE",X"C2",X"C3",X"C7",X"C4",X"C5",X"C0",X"FF",X"10",X"C9",
		X"CE",X"CA",X"CB",X"CF",X"CC",X"CD",X"A0",X"FF",X"D8",X"D9",X"DA",X"DB",X"DC",X"DD",X"DE",X"DF",
		X"3E",X"C8",X"3E",X"C8",X"74",X"54",X"74",X"54",X"3A",X"30",X"8F",X"E6",X"07",X"EF",X"8F",X"27",
		X"F3",X"27",X"56",X"28",X"AD",X"28",X"C5",X"28",X"26",X"80",X"77",X"D7",X"0D",X"20",X"FA",X"3A",
		X"3F",X"8F",X"A7",X"20",X"1D",X"3A",X"75",X"8D",X"A7",X"28",X"0A",X"21",X"20",X"8F",X"7E",X"A7",
		X"20",X"03",X"34",X"18",X"08",X"3A",X"01",X"89",X"A7",X"C8",X"E6",X"07",X"C0",X"3E",X"01",X"32",
		X"3F",X"8F",X"3A",X"B4",X"8A",X"FE",X"3C",X"D8",X"3A",X"90",X"8C",X"CB",X"4F",X"C0",X"3A",X"A8",
		X"8C",X"CB",X"4F",X"C0",X"21",X"30",X"8F",X"34",X"3E",X"08",X"32",X"2F",X"89",X"3A",X"06",X"88",
		X"A7",X"20",X"0E",X"3A",X"50",X"8F",X"21",X"3F",X"8F",X"B6",X"28",X"05",X"3E",X"6F",X"32",X"08",
		X"85",X"3A",X"7A",X"8D",X"A7",X"28",X"03",X"32",X"20",X"8F",X"21",X"A7",X"84",X"11",X"51",X"2D",
		X"C3",X"25",X"33",X"3A",X"B4",X"8A",X"FE",X"34",X"38",X"19",X"21",X"2F",X"89",X"35",X"C0",X"36",
		X"10",X"2B",X"34",X"CB",X"46",X"21",X"A7",X"84",X"11",X"51",X"2D",X"20",X"03",X"11",X"55",X"2D",
		X"C3",X"25",X"33",X"21",X"90",X"8C",X"11",X"18",X"00",X"06",X"02",X"7E",X"A7",X"28",X"04",X"19",
		X"10",X"F9",X"C9",X"3E",X"02",X"32",X"30",X"8F",X"77",X"CD",X"05",X"0F",X"21",X"A7",X"84",X"11",
		X"55",X"2D",X"CD",X"25",X"33",X"3A",X"50",X"8F",X"21",X"3F",X"8F",X"B6",X"28",X"03",X"3E",X"10",
		X"32",X"08",X"85",X"3E",X"01",X"32",X"99",X"8A",X"3A",X"86",X"8A",X"C6",X"0C",X"32",X"9E",X"8A",
		X"3E",X"10",X"32",X"A7",X"8A",X"C9",X"3A",X"50",X"8F",X"A7",X"20",X"3A",X"DD",X"21",X"78",X"8C",
		X"11",X"E8",X"FF",X"06",X"06",X"DD",X"7E",X"00",X"DD",X"B6",X"01",X"28",X"05",X"DD",X"19",X"10",
		X"F4",X"C9",X"DD",X"36",X"01",X"05",X"DD",X"36",X"02",X"10",X"DD",X"36",X"03",X"00",X"DD",X"36",
		X"04",X"08",X"DD",X"36",X"05",X"00",X"DD",X"36",X"06",X"1A",X"DD",X"36",X"0F",X"37",X"DD",X"36",
		X"10",X"42",X"DD",X"22",X"32",X"8F",X"21",X"30",X"8F",X"34",X"3A",X"61",X"8F",X"A7",X"28",X"04",
		X"2E",X"5D",X"34",X"C9",X"2E",X"34",X"36",X"20",X"11",X"15",X"03",X"FF",X"C9",X"21",X"34",X"8F",
		X"7E",X"A7",X"28",X"02",X"35",X"C9",X"2E",X"30",X"34",X"3A",X"50",X"8F",X"A7",X"C0",X"AF",X"2A",
		X"32",X"8F",X"06",X"18",X"D7",X"C9",X"CD",X"01",X"21",X"3A",X"07",X"89",X"CB",X"47",X"21",X"0A",
		X"88",X"20",X"03",X"36",X"06",X"C9",X"3A",X"08",X"8F",X"A7",X"28",X"03",X"36",X"04",X"C9",X"DD",
		X"21",X"80",X"8A",X"21",X"8D",X"2B",X"E5",X"DD",X"35",X"11",X"C0",X"DD",X"7E",X"02",X"E6",X"07",
		X"EF",X"01",X"29",X"A0",X"29",X"01",X"2A",X"32",X"2A",X"79",X"2A",X"96",X"2A",X"B3",X"2A",X"E8",
		X"2A",X"DD",X"36",X"11",X"01",X"DD",X"34",X"04",X"DD",X"7E",X"04",X"FE",X"DC",X"30",X"0F",X"CD",
		X"D7",X"23",X"3A",X"BE",X"88",X"FE",X"F9",X"C8",X"CD",X"05",X"24",X"C3",X"A1",X"23",X"21",X"59",
		X"2D",X"CD",X"0F",X"25",X"21",X"91",X"8A",X"36",X"0C",X"2E",X"82",X"34",X"23",X"23",X"7E",X"D6",
		X"03",X"77",X"AF",X"32",X"9C",X"8A",X"32",X"9E",X"8A",X"21",X"59",X"08",X"01",X"00",X"20",X"7E",
		X"81",X"4F",X"23",X"10",X"FA",X"FE",X"63",X"C2",X"E8",X"2A",X"06",X"20",X"11",X"80",X"29",X"1B",
		X"1A",X"BE",X"C2",X"9A",X"2B",X"23",X"10",X"F7",X"CD",X"A2",X"0F",X"C9",X"D2",X"24",X"30",X"14",
		X"11",X"10",X"10",X"12",X"12",X"12",X"12",X"12",X"12",X"12",X"12",X"12",X"12",X"12",X"12",X"12",
		X"12",X"12",X"12",X"12",X"12",X"12",X"12",X"12",X"12",X"12",X"12",X"12",X"12",X"12",X"03",X"1D",
		X"0D",X"03",X"00",X"00",X"07",X"07",X"07",X"07",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0B",X"0B",X"0B",X"0B",X"07",X"00",X"04",X"00",
		X"DD",X"36",X"11",X"03",X"DD",X"34",X"0B",X"DD",X"7E",X"0B",X"E6",X"03",X"20",X"0E",X"DD",X"7E",
		X"0F",X"FE",X"15",X"3E",X"15",X"20",X"02",X"3E",X"1E",X"DD",X"77",X"0F",X"DD",X"7E",X"06",X"D6",
		X"02",X"DD",X"77",X"06",X"FE",X"2C",X"D0",X"3A",X"43",X"83",X"A7",X"C2",X"23",X"2B",X"C6",X"30",
		X"32",X"30",X"8D",X"DD",X"36",X"11",X"18",X"DD",X"34",X"02",X"21",X"79",X"08",X"01",X"00",X"20",
		X"7E",X"81",X"4F",X"23",X"10",X"FA",X"FE",X"37",X"C2",X"B3",X"2A",X"21",X"59",X"08",X"06",X"20",
		X"11",X"80",X"29",X"1A",X"BE",X"C2",X"01",X"29",X"23",X"13",X"10",X"F7",X"11",X"14",X"06",X"FF",
		X"C9",X"DD",X"36",X"11",X"08",X"DD",X"CB",X"10",X"FE",X"21",X"5A",X"87",X"3E",X"BC",X"77",X"23",
		X"77",X"23",X"77",X"DD",X"34",X"02",X"AF",X"21",X"39",X"08",X"06",X"20",X"86",X"23",X"10",X"FC",
		X"3D",X"C2",X"58",X"2C",X"11",X"15",X"06",X"FF",X"21",X"03",X"89",X"7E",X"FE",X"09",X"D8",X"36",
		X"08",X"C9",X"DD",X"36",X"11",X"03",X"DD",X"34",X"0B",X"DD",X"7E",X"0B",X"E6",X"03",X"20",X"0E",
		X"DD",X"7E",X"0F",X"FE",X"15",X"3E",X"15",X"20",X"02",X"3E",X"1E",X"DD",X"77",X"0F",X"3E",X"80",
		X"DD",X"86",X"05",X"DD",X"77",X"05",X"DD",X"7E",X"06",X"30",X"01",X"3C",X"3C",X"DD",X"77",X"06",
		X"FE",X"52",X"20",X"05",X"11",X"94",X"06",X"FF",X"C9",X"FE",X"64",X"20",X"05",X"11",X"95",X"06",
		X"FF",X"C9",X"FE",X"AC",X"D8",X"DD",X"34",X"02",X"C9",X"21",X"66",X"1C",X"11",X"23",X"2B",X"06",
		X"68",X"1A",X"96",X"C2",X"A0",X"29",X"23",X"13",X"10",X"F7",X"DD",X"36",X"11",X"30",X"DD",X"CB",
		X"10",X"BE",X"DD",X"34",X"02",X"C9",X"21",X"DF",X"67",X"11",X"23",X"2B",X"06",X"20",X"1A",X"96",
		X"C2",X"01",X"2A",X"23",X"1B",X"10",X"F7",X"DD",X"36",X"11",X"18",X"DD",X"CB",X"10",X"FE",X"DD",
		X"34",X"02",X"C9",X"DD",X"36",X"11",X"02",X"DD",X"34",X"0B",X"DD",X"7E",X"0B",X"E6",X"03",X"20",
		X"0E",X"DD",X"7E",X"0F",X"FE",X"15",X"3E",X"15",X"20",X"02",X"3E",X"1E",X"DD",X"77",X"0F",X"DD",
		X"34",X"06",X"DD",X"7E",X"06",X"FE",X"C0",X"D8",X"DD",X"7E",X"04",X"D6",X"03",X"DD",X"77",X"04",
		X"DD",X"34",X"02",X"DD",X"36",X"11",X"40",X"C9",X"AF",X"21",X"80",X"8A",X"77",X"11",X"81",X"8A",
		X"01",X"40",X"02",X"ED",X"B0",X"32",X"02",X"89",X"32",X"03",X"89",X"32",X"31",X"89",X"3E",X"06",
		X"32",X"0A",X"88",X"C9",X"AF",X"88",X"0A",X"32",X"88",X"08",X"32",X"89",X"04",X"32",X"01",X"3E",
		X"AD",X"20",X"B9",X"5A",X"3E",X"FA",X"10",X"19",X"4F",X"81",X"7E",X"0A",X"00",X"01",X"FF",X"E0",
		X"11",X"82",X"BC",X"21",X"08",X"88",X"35",X"3A",X"2A",X"8E",X"A7",X"28",X"04",X"7E",X"A7",X"28",
		X"28",X"CD",X"94",X"7E",X"3A",X"FC",X"89",X"A7",X"C8",X"3A",X"08",X"88",X"E6",X"07",X"C0",X"3A",
		X"FF",X"89",X"2A",X"FD",X"89",X"11",X"20",X"00",X"06",X"1C",X"77",X"19",X"10",X"FC",X"3C",X"FE",
		X"10",X"38",X"02",X"3E",X"06",X"32",X"FF",X"89",X"C9",X"21",X"5F",X"85",X"11",X"E0",X"FF",X"06",
		X"08",X"3E",X"10",X"77",X"19",X"10",X"FA",X"21",X"BC",X"82",X"11",X"E0",X"FF",X"01",X"00",X"0A",
		X"7E",X"81",X"4F",X"19",X"10",X"FA",X"79",X"FE",X"AA",X"C0",X"AF",X"32",X"2A",X"8E",X"3A",X"0E",
		X"88",X"A7",X"28",X"4E",X"3A",X"0D",X"88",X"A7",X"28",X"29",X"3A",X"48",X"89",X"3A",X"82",X"8A",
		X"FE",X"03",X"D8",X"CD",X"9A",X"2B",X"CD",X"2C",X"2C",X"C9",X"21",X"03",X"89",X"7E",X"FE",X"02",
		X"DC",X"BF",X"2B",X"21",X"30",X"8D",X"7E",X"A7",X"28",X"02",X"35",X"C9",X"DD",X"21",X"60",X"8C",
		X"11",X"E8",X"FF",X"06",X"11",X"D9",X"CD",X"E5",X"2B",X"D9",X"DD",X"19",X"10",X"F7",X"C9",X"FE",
		X"01",X"21",X"7B",X"87",X"28",X"0D",X"7E",X"FE",X"BA",X"20",X"02",X"F1",X"C9",X"11",X"E1",X"2B",
		X"CD",X"25",X"33",X"21",X"BB",X"87",X"7E",X"FE",X"BA",X"C8",X"11",X"E1",X"2B",X"CD",X"25",X"33",
		X"C9",X"BA",X"BA",X"BA",X"BA",X"DD",X"7E",X"00",X"DD",X"B6",X"01",X"0F",X"D8",X"DD",X"36",X"00",
		X"01",X"AF",X"DD",X"36",X"02",X"11",X"DD",X"77",X"03",X"DD",X"77",X"05",X"DD",X"36",X"04",X"1C",
		X"DD",X"36",X"06",X"03",X"21",X"03",X"89",X"35",X"CB",X"46",X"28",X"01",X"3C",X"DD",X"77",X"07",
		X"11",X"5D",X"2D",X"CD",X"1E",X"38",X"3A",X"03",X"89",X"FE",X"0A",X"38",X"02",X"3E",X"0A",X"47",
		X"3E",X"20",X"90",X"32",X"30",X"8D",X"DD",X"36",X"09",X"10",X"F1",X"C9",X"DD",X"21",X"E0",X"8A",
		X"11",X"18",X"00",X"06",X"11",X"D9",X"CD",X"3F",X"2C",X"D9",X"DD",X"19",X"10",X"F7",X"C9",X"DD",
		X"7E",X"00",X"DD",X"B6",X"01",X"0F",X"D0",X"DD",X"7E",X"02",X"E6",X"1F",X"D6",X"11",X"D8",X"EF",
		X"58",X"2C",X"B3",X"2C",X"24",X"2D",X"4A",X"2D",X"CD",X"06",X"40",X"DD",X"7E",X"05",X"DD",X"86",
		X"09",X"30",X"03",X"DD",X"34",X"06",X"DD",X"77",X"05",X"47",X"DD",X"7E",X"06",X"FE",X"12",X"D8",
		X"DD",X"21",X"E0",X"8A",X"06",X"11",X"CD",X"85",X"2C",X"11",X"18",X"00",X"DD",X"19",X"10",X"F6",
		X"CD",X"3F",X"0F",X"F1",X"C9",X"DD",X"7E",X"02",X"FE",X"11",X"C0",X"DD",X"36",X"02",X"12",X"11",
		X"A7",X"2C",X"CD",X"1E",X"38",X"21",X"00",X"2D",X"DD",X"75",X"16",X"DD",X"74",X"17",X"DD",X"36",
		X"15",X"00",X"C9",X"A7",X"2C",X"AD",X"2C",X"4F",X"04",X"F0",X"FF",X"A7",X"2C",X"0F",X"04",X"F0",
		X"FF",X"AD",X"2C",X"CD",X"06",X"40",X"DD",X"6E",X"16",X"DD",X"66",X"17",X"7E",X"FE",X"FF",X"20",
		X"06",X"DD",X"77",X"15",X"23",X"18",X"F5",X"FE",X"88",X"20",X"0E",X"DD",X"34",X"02",X"11",X"5D",
		X"2D",X"CD",X"1E",X"38",X"DD",X"36",X"11",X"20",X"C9",X"23",X"DD",X"75",X"16",X"DD",X"74",X"17",
		X"DD",X"CB",X"15",X"46",X"20",X"0E",X"47",X"DD",X"7E",X"03",X"90",X"30",X"03",X"DD",X"35",X"04",
		X"DD",X"77",X"03",X"C9",X"DD",X"86",X"03",X"30",X"03",X"DD",X"34",X"04",X"DD",X"77",X"03",X"C9",
		X"C0",X"80",X"60",X"40",X"40",X"20",X"20",X"20",X"00",X"20",X"00",X"20",X"00",X"00",X"20",X"00",
		X"00",X"FF",X"00",X"00",X"20",X"00",X"00",X"20",X"00",X"20",X"00",X"20",X"20",X"20",X"40",X"40",
		X"60",X"80",X"C0",X"88",X"CD",X"06",X"40",X"DD",X"7E",X"05",X"DD",X"86",X"09",X"30",X"03",X"DD",
		X"34",X"06",X"DD",X"77",X"05",X"DD",X"7E",X"06",X"FE",X"19",X"D8",X"DD",X"34",X"02",X"AF",X"DD",
		X"77",X"05",X"DD",X"77",X"06",X"DD",X"77",X"16",X"F1",X"C9",X"3E",X"00",X"32",X"36",X"8F",X"F1",
		X"C9",X"F0",X"F1",X"F3",X"F2",X"A2",X"A1",X"10",X"10",X"15",X"00",X"0A",X"0F",X"40",X"03",X"07",
		X"40",X"09",X"07",X"FF",X"5D",X"2D",X"3A",X"32",X"8D",X"A7",X"C0",X"3A",X"03",X"89",X"D6",X"02",
		X"C8",X"CD",X"78",X"2D",X"CD",X"22",X"2E",X"C9",X"3A",X"14",X"8F",X"EF",X"80",X"2D",X"BC",X"2D",
		X"3A",X"03",X"89",X"D6",X"02",X"21",X"31",X"89",X"BE",X"C8",X"34",X"21",X"18",X"8F",X"7E",X"FE",
		X"04",X"38",X"05",X"3A",X"EF",X"89",X"A7",X"C8",X"34",X"21",X"B8",X"2D",X"E7",X"6F",X"26",X"84",
		X"22",X"19",X"8F",X"3A",X"18",X"8F",X"47",X"21",X"26",X"8F",X"23",X"23",X"10",X"FC",X"36",X"10",
		X"2E",X"14",X"34",X"2E",X"16",X"36",X"10",X"C9",X"97",X"93",X"8F",X"8A",X"21",X"16",X"8F",X"7E",
		X"A7",X"28",X"02",X"35",X"C9",X"36",X"08",X"2E",X"1B",X"7E",X"FE",X"08",X"20",X"0F",X"AF",X"77",
		X"2E",X"14",X"77",X"3A",X"18",X"8F",X"2E",X"1B",X"85",X"6F",X"36",X"01",X"C9",X"21",X"EE",X"2D",
		X"CD",X"45",X"0C",X"2A",X"19",X"8F",X"CD",X"25",X"33",X"21",X"1B",X"8F",X"34",X"C9",X"FE",X"2D",
		X"02",X"2E",X"06",X"2E",X"0A",X"2E",X"0E",X"2E",X"12",X"2E",X"16",X"2E",X"1A",X"2E",X"39",X"39",
		X"3A",X"3A",X"39",X"F4",X"F6",X"3A",X"39",X"F5",X"F7",X"3A",X"39",X"F8",X"FA",X"3A",X"F4",X"FC",
		X"FE",X"F6",X"F5",X"FD",X"FF",X"F7",X"F8",X"E0",X"E2",X"FA",X"F9",X"E1",X"E3",X"FB",X"39",X"39",
		X"A7",X"A6",X"3A",X"18",X"8F",X"A7",X"C8",X"DD",X"21",X"1C",X"8F",X"47",X"D9",X"CD",X"36",X"2E",
		X"D9",X"DD",X"23",X"10",X"F7",X"C9",X"DD",X"7E",X"00",X"D6",X"01",X"D8",X"EF",X"5E",X"2E",X"CB",
		X"2E",X"01",X"2F",X"2F",X"2F",X"DD",X"7D",X"4F",X"E6",X"03",X"87",X"C6",X"28",X"6F",X"26",X"8F",
		X"35",X"C9",X"DD",X"7D",X"E6",X"03",X"21",X"B8",X"2D",X"E7",X"6F",X"26",X"84",X"C9",X"3A",X"5F",
		X"8A",X"E6",X"03",X"C0",X"CD",X"45",X"2E",X"C0",X"36",X"01",X"FD",X"21",X"48",X"8C",X"11",X"18",
		X"00",X"06",X"03",X"FD",X"7E",X"00",X"FD",X"B6",X"01",X"0F",X"30",X"05",X"FD",X"19",X"10",X"F3",
		X"C9",X"3A",X"07",X"89",X"FE",X"10",X"38",X"02",X"3E",X"10",X"D6",X"28",X"2F",X"77",X"23",X"78",
		X"2F",X"E6",X"03",X"77",X"DD",X"7D",X"E6",X"03",X"21",X"C7",X"2E",X"E7",X"FD",X"36",X"00",X"07",
		X"FD",X"36",X"02",X"10",X"FD",X"77",X"04",X"FD",X"36",X"05",X"40",X"FD",X"36",X"06",X"1A",X"FD",
		X"36",X"0F",X"2E",X"FD",X"36",X"10",X"40",X"DD",X"34",X"00",X"CD",X"52",X"2E",X"11",X"FE",X"2D",
		X"CD",X"25",X"33",X"CD",X"11",X"0F",X"C9",X"18",X"14",X"10",X"0B",X"CD",X"45",X"2E",X"C0",X"3A",
		X"07",X"89",X"FE",X"10",X"38",X"02",X"3E",X"10",X"07",X"C6",X"18",X"77",X"FD",X"21",X"30",X"8C",
		X"11",X"18",X"00",X"23",X"46",X"04",X"FD",X"19",X"10",X"FC",X"FD",X"34",X"0F",X"FD",X"36",X"05",
		X"00",X"FD",X"35",X"06",X"DD",X"34",X"00",X"CD",X"52",X"2E",X"11",X"1E",X"2E",X"CD",X"25",X"33",
		X"C9",X"CD",X"5F",X"30",X"CD",X"45",X"2E",X"C0",X"36",X"0C",X"FD",X"21",X"30",X"8C",X"11",X"18",
		X"00",X"23",X"46",X"04",X"FD",X"19",X"10",X"FC",X"FD",X"35",X"0F",X"FD",X"36",X"05",X"C0",X"FD",
		X"34",X"06",X"DD",X"34",X"00",X"CD",X"52",X"2E",X"11",X"FE",X"2D",X"CD",X"25",X"33",X"C9",X"CD",
		X"45",X"2E",X"C0",X"3A",X"31",X"89",X"A7",X"C8",X"E5",X"3A",X"07",X"89",X"CB",X"3F",X"CB",X"3F",
		X"FE",X"04",X"38",X"02",X"3E",X"03",X"47",X"3A",X"20",X"88",X"E6",X"04",X"0F",X"80",X"21",X"93",
		X"2F",X"CD",X"45",X"0C",X"EB",X"3A",X"31",X"89",X"3D",X"FE",X"20",X"38",X"02",X"3E",X"1F",X"E7",
		X"E1",X"5F",X"7D",X"FE",X"28",X"28",X"0C",X"D6",X"02",X"6F",X"7E",X"E6",X"1C",X"83",X"5F",X"7D",
		X"C6",X"02",X"6F",X"7B",X"77",X"11",X"18",X"00",X"23",X"46",X"21",X"30",X"8C",X"04",X"19",X"10",
		X"FD",X"AF",X"06",X"18",X"D7",X"3C",X"DD",X"77",X"00",X"CD",X"52",X"2E",X"11",X"1A",X"2E",X"CD",
		X"25",X"33",X"C9",X"9F",X"2F",X"BF",X"2F",X"DF",X"2F",X"FF",X"2F",X"1F",X"30",X"3F",X"30",X"64",
		X"64",X"60",X"60",X"60",X"5C",X"5C",X"58",X"58",X"58",X"4C",X"4C",X"48",X"48",X"48",X"40",X"40",
		X"40",X"3C",X"3C",X"3C",X"38",X"38",X"30",X"30",X"30",X"2C",X"2C",X"20",X"20",X"18",X"10",X"58",
		X"58",X"58",X"54",X"54",X"50",X"50",X"4C",X"4C",X"48",X"48",X"40",X"40",X"40",X"3C",X"3C",X"38",
		X"38",X"34",X"34",X"30",X"30",X"2C",X"2C",X"28",X"28",X"24",X"24",X"18",X"18",X"10",X"08",X"48",
		X"48",X"48",X"44",X"3C",X"3C",X"34",X"34",X"30",X"30",X"28",X"28",X"24",X"24",X"20",X"20",X"1C",
		X"1C",X"18",X"18",X"14",X"14",X"10",X"10",X"0C",X"0C",X"08",X"08",X"04",X"04",X"03",X"02",X"38",
		X"38",X"34",X"34",X"2C",X"2C",X"28",X"28",X"24",X"24",X"20",X"20",X"1C",X"1C",X"18",X"18",X"14",
		X"14",X"10",X"10",X"0C",X"0C",X"08",X"08",X"04",X"04",X"04",X"04",X"02",X"02",X"02",X"01",X"20",
		X"20",X"20",X"1C",X"1C",X"18",X"18",X"14",X"14",X"10",X"10",X"10",X"0C",X"0C",X"0C",X"08",X"08",
		X"08",X"04",X"04",X"04",X"02",X"02",X"02",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"18",
		X"18",X"18",X"18",X"14",X"14",X"14",X"10",X"10",X"10",X"0C",X"0C",X"0C",X"08",X"08",X"04",X"04",
		X"04",X"02",X"02",X"02",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"DD",
		X"7D",X"E6",X"03",X"21",X"87",X"30",X"E7",X"47",X"3A",X"84",X"8A",X"D6",X"07",X"4F",X"C6",X"0E",
		X"B8",X"D8",X"79",X"B8",X"D0",X"21",X"24",X"8F",X"3A",X"08",X"8F",X"B6",X"C0",X"3E",X"01",X"32",
		X"32",X"8D",X"CD",X"15",X"0F",X"F1",X"C9",X"C0",X"A0",X"80",X"58",X"3A",X"04",X"8F",X"A7",X"C8",
		X"3A",X"08",X"8F",X"A7",X"20",X"4A",X"DD",X"21",X"E0",X"8A",X"FD",X"21",X"20",X"89",X"11",X"18",
		X"00",X"06",X"11",X"DD",X"7E",X"00",X"A7",X"28",X"0D",X"FE",X"05",X"28",X"09",X"DD",X"19",X"10",
		X"F2",X"AF",X"32",X"20",X"89",X"C9",X"DD",X"7E",X"01",X"A7",X"20",X"F1",X"DD",X"E5",X"E1",X"FD",
		X"75",X"00",X"FD",X"74",X"01",X"DD",X"36",X"00",X"05",X"DD",X"36",X"02",X"10",X"FD",X"23",X"FD",
		X"23",X"FD",X"7D",X"FE",X"28",X"20",X"D6",X"21",X"08",X"8F",X"36",X"01",X"23",X"36",X"20",X"C9",
		X"21",X"BD",X"32",X"E5",X"3A",X"08",X"8F",X"E6",X"03",X"3D",X"EF",X"F1",X"30",X"6E",X"31",X"66",
		X"32",X"DD",X"21",X"20",X"89",X"21",X"37",X"33",X"06",X"04",X"DD",X"5E",X"00",X"DD",X"56",X"01",
		X"FD",X"6B",X"FD",X"62",X"7E",X"FD",X"77",X"04",X"23",X"7E",X"FD",X"77",X"06",X"23",X"7E",X"FD",
		X"77",X"0F",X"23",X"7E",X"FD",X"77",X"10",X"FD",X"36",X"09",X"30",X"DD",X"23",X"DD",X"23",X"23",
		X"10",X"D8",X"3E",X"0C",X"32",X"28",X"89",X"21",X"08",X"8F",X"34",X"3E",X"10",X"11",X"1D",X"00",
		X"21",X"C2",X"84",X"0E",X"03",X"06",X"03",X"D7",X"19",X"0D",X"20",X"F9",X"21",X"70",X"33",X"22",
		X"4B",X"8F",X"CD",X"19",X"0F",X"CD",X"3E",X"32",X"11",X"AC",X"68",X"21",X"78",X"32",X"06",X"40",
		X"7B",X"BE",X"20",X"0F",X"7A",X"23",X"BE",X"20",X"0A",X"23",X"1A",X"BE",X"20",X"05",X"13",X"23",
		X"10",X"F8",X"C9",X"AF",X"21",X"00",X"88",X"11",X"01",X"88",X"77",X"ED",X"B0",X"C9",X"21",X"28",
		X"89",X"7E",X"A7",X"28",X"02",X"35",X"C9",X"2E",X"20",X"5E",X"23",X"56",X"D5",X"FD",X"E1",X"2A",
		X"4B",X"8F",X"7E",X"A7",X"28",X"13",X"FD",X"86",X"05",X"30",X"03",X"FD",X"34",X"06",X"FD",X"77",
		X"05",X"23",X"7E",X"23",X"22",X"4B",X"8F",X"18",X"0B",X"FD",X"34",X"09",X"20",X"03",X"FD",X"34",
		X"04",X"FD",X"7E",X"09",X"FD",X"86",X"03",X"30",X"03",X"FD",X"34",X"04",X"FD",X"77",X"03",X"3A",
		X"4A",X"8F",X"A7",X"FD",X"7E",X"04",X"20",X"1F",X"07",X"07",X"07",X"C6",X"18",X"4F",X"3A",X"84",
		X"8A",X"B9",X"30",X"21",X"3E",X"01",X"32",X"24",X"8F",X"32",X"4A",X"8F",X"21",X"48",X"33",X"22",
		X"4B",X"8F",X"CD",X"1D",X"0F",X"18",X"0E",X"FE",X"1B",X"38",X"0A",X"32",X"28",X"89",X"21",X"08",
		X"8F",X"34",X"CD",X"1D",X"0F",X"FD",X"4E",X"04",X"FD",X"46",X"06",X"DD",X"21",X"20",X"89",X"11",
		X"03",X"00",X"DD",X"6E",X"02",X"DD",X"66",X"03",X"19",X"FD",X"7E",X"03",X"77",X"23",X"79",X"77",
		X"23",X"FD",X"7E",X"05",X"77",X"23",X"78",X"C6",X"02",X"77",X"DD",X"6E",X"04",X"DD",X"66",X"05",
		X"19",X"FD",X"7E",X"03",X"77",X"23",X"79",X"C6",X"02",X"77",X"23",X"FD",X"7E",X"05",X"77",X"23",
		X"78",X"77",X"DD",X"6E",X"06",X"DD",X"66",X"07",X"19",X"FD",X"7E",X"03",X"77",X"23",X"79",X"C6",
		X"02",X"77",X"23",X"FD",X"7E",X"05",X"77",X"23",X"78",X"C6",X"02",X"77",X"06",X"04",X"DD",X"7E",
		X"01",X"FE",X"8C",X"CC",X"4D",X"32",X"DD",X"23",X"DD",X"23",X"10",X"F2",X"C9",X"DD",X"7E",X"00",
		X"FE",X"40",X"D8",X"26",X"8C",X"C6",X"05",X"6F",X"7E",X"D6",X"40",X"77",X"D0",X"23",X"35",X"3A",
		X"E5",X"89",X"A7",X"20",X"13",X"C9",X"21",X"99",X"07",X"01",X"00",X"20",X"7E",X"81",X"4F",X"23",
		X"10",X"FA",X"FE",X"DC",X"C2",X"99",X"07",X"C9",X"AC",X"68",X"21",X"55",X"8F",X"7E",X"A7",X"C0",
		X"34",X"21",X"02",X"84",X"11",X"00",X"00",X"7E",X"83",X"5F",X"30",X"01",X"14",X"2C",X"7D",X"E6",
		X"1F",X"FE",X"1F",X"20",X"F2",X"7D",X"C6",X"03",X"6F",X"30",X"EC",X"24",X"7C",X"FE",X"88",X"38",
		X"E6",X"21",X"EB",X"68",X"06",X"04",X"7B",X"BE",X"28",X"06",X"23",X"10",X"FA",X"C3",X"D4",X"76",
		X"7A",X"23",X"BE",X"C8",X"10",X"FA",X"C3",X"29",X"38",X"43",X"95",X"89",X"87",X"3A",X"24",X"8F",
		X"A7",X"C8",X"FE",X"02",X"28",X"22",X"D0",X"AF",X"21",X"21",X"8D",X"77",X"23",X"36",X"20",X"CD",
		X"AD",X"0F",X"21",X"24",X"8F",X"34",X"21",X"79",X"07",X"01",X"00",X"20",X"7E",X"81",X"4F",X"23",
		X"10",X"FA",X"E6",X"47",X"C2",X"40",X"1F",X"C9",X"21",X"84",X"8A",X"34",X"34",X"7E",X"FE",X"DB",
		X"30",X"04",X"CD",X"D7",X"23",X"C9",X"CD",X"30",X"0F",X"3A",X"83",X"80",X"A7",X"C0",X"3C",X"32",
		X"32",X"8D",X"21",X"24",X"8F",X"34",X"C9",X"01",X"1D",X"00",X"C5",X"06",X"03",X"1A",X"77",X"13",
		X"23",X"10",X"FA",X"C1",X"09",X"3A",X"0B",X"8F",X"3C",X"32",X"0B",X"8F",X"FE",X"03",X"20",X"E7",
		X"AF",X"32",X"0B",X"8F",X"C9",X"01",X"20",X"00",X"1A",X"77",X"13",X"23",X"1A",X"77",X"13",X"09",
		X"1A",X"77",X"13",X"2B",X"1A",X"77",X"C9",X"02",X"17",X"30",X"40",X"02",X"19",X"35",X"40",X"04",
		X"17",X"38",X"40",X"04",X"19",X"3F",X"40",X"FF",X"20",X"00",X"20",X"00",X"20",X"00",X"20",X"00",
		X"20",X"10",X"20",X"10",X"20",X"10",X"20",X"10",X"20",X"18",X"20",X"18",X"20",X"18",X"20",X"18",
		X"18",X"20",X"18",X"20",X"18",X"20",X"18",X"20",X"10",X"28",X"10",X"28",X"10",X"28",X"10",X"28",
		X"10",X"30",X"10",X"30",X"10",X"30",X"00",X"DD",X"21",X"E0",X"8A",X"11",X"18",X"00",X"06",X"0E",
		X"D9",X"CD",X"8A",X"33",X"D9",X"DD",X"19",X"10",X"F7",X"C9",X"DD",X"7E",X"00",X"DD",X"B6",X"01",
		X"0F",X"D0",X"DD",X"7E",X"02",X"E6",X"1F",X"FE",X"11",X"D0",X"EF",X"BD",X"33",X"23",X"34",X"36",
		X"35",X"5B",X"35",X"65",X"38",X"AF",X"39",X"E3",X"3B",X"92",X"3C",X"18",X"3D",X"5C",X"3D",X"8F",
		X"3D",X"69",X"3E",X"9C",X"3E",X"5C",X"3F",X"72",X"3F",X"7C",X"3F",X"E9",X"3F",X"DD",X"35",X"11",
		X"C0",X"DD",X"34",X"02",X"DD",X"CB",X"0B",X"46",X"20",X"2D",X"3A",X"43",X"8D",X"E6",X"0F",X"21",
		X"18",X"34",X"E7",X"32",X"4B",X"8D",X"DD",X"BE",X"06",X"28",X"11",X"3E",X"00",X"11",X"29",X"38",
		X"30",X"04",X"3C",X"11",X"38",X"38",X"DD",X"77",X"08",X"C3",X"1E",X"38",X"DD",X"7E",X"09",X"DD",
		X"BE",X"05",X"38",X"EF",X"C3",X"73",X"34",X"21",X"4C",X"8D",X"34",X"3E",X"06",X"32",X"01",X"89",
		X"AF",X"32",X"4A",X"8D",X"DD",X"77",X"0B",X"CD",X"CA",X"33",X"11",X"47",X"38",X"DD",X"CB",X"08",
		X"46",X"28",X"D6",X"11",X"56",X"38",X"18",X"D1",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"00",
		X"00",X"00",X"00",X"CD",X"06",X"40",X"DD",X"CB",X"01",X"46",X"28",X"0B",X"3A",X"63",X"8F",X"A7",
		X"C0",X"DD",X"36",X"01",X"00",X"18",X"3C",X"DD",X"7E",X"08",X"A7",X"C2",X"F2",X"34",X"DD",X"7E",
		X"05",X"DD",X"86",X"09",X"30",X"03",X"DD",X"34",X"06",X"DD",X"77",X"05",X"47",X"3A",X"4B",X"8D",
		X"4F",X"DD",X"7E",X"06",X"E6",X"1F",X"B9",X"D8",X"28",X"0A",X"DD",X"36",X"08",X"01",X"11",X"38",
		X"38",X"C3",X"1E",X"38",X"A7",X"CA",X"B0",X"34",X"3A",X"0A",X"88",X"FE",X"04",X"C0",X"DD",X"7E",
		X"09",X"B8",X"D8",X"3A",X"63",X"8F",X"A7",X"CA",X"7F",X"34",X"DD",X"36",X"01",X"01",X"C9",X"DD",
		X"36",X"01",X"00",X"21",X"43",X"8D",X"7E",X"FE",X"07",X"30",X"25",X"FE",X"0A",X"30",X"01",X"34",
		X"7E",X"21",X"18",X"34",X"E7",X"32",X"4B",X"8D",X"21",X"E3",X"86",X"11",X"40",X"00",X"36",X"D8",
		X"23",X"36",X"D9",X"1E",X"1F",X"19",X"36",X"DA",X"23",X"36",X"DB",X"3E",X"01",X"32",X"63",X"8F",
		X"CD",X"53",X"35",X"21",X"40",X"8D",X"35",X"21",X"01",X"89",X"7E",X"4F",X"A7",X"28",X"01",X"35",
		X"3A",X"0A",X"88",X"FE",X"04",X"20",X"02",X"2C",X"34",X"3A",X"01",X"89",X"47",X"21",X"43",X"87",
		X"11",X"20",X"00",X"FE",X"0A",X"38",X"0C",X"3A",X"50",X"8F",X"A7",X"C0",X"AF",X"C6",X"01",X"27",
		X"10",X"FB",X"47",X"E6",X"0F",X"77",X"19",X"78",X"0F",X"0F",X"0F",X"0F",X"E6",X"0F",X"A7",X"C8",
		X"77",X"C9",X"DD",X"7E",X"0A",X"ED",X"44",X"47",X"DD",X"7E",X"05",X"B8",X"30",X"03",X"DD",X"35",
		X"06",X"DD",X"86",X"0A",X"DD",X"77",X"05",X"47",X"3A",X"4B",X"8D",X"4F",X"DD",X"7E",X"06",X"E6",
		X"1F",X"B9",X"28",X"10",X"D0",X"A7",X"CA",X"B0",X"34",X"3A",X"0A",X"88",X"FE",X"04",X"C0",X"DD",
		X"36",X"08",X"00",X"C9",X"A7",X"CA",X"B0",X"34",X"3A",X"0A",X"88",X"FE",X"04",X"C0",X"DD",X"7E",
		X"09",X"B8",X"D8",X"C3",X"73",X"34",X"CD",X"06",X"40",X"DD",X"35",X"11",X"C0",X"DD",X"7E",X"07",
		X"E6",X"F0",X"28",X"0F",X"21",X"76",X"8D",X"34",X"7E",X"FE",X"03",X"38",X"06",X"2D",X"AF",X"77",
		X"32",X"20",X"8F",X"AF",X"DD",X"E5",X"E1",X"06",X"17",X"D7",X"C9",X"CD",X"06",X"40",X"DD",X"7E",
		X"08",X"A7",X"C2",X"57",X"37",X"DD",X"7E",X"05",X"DD",X"86",X"09",X"30",X"03",X"DD",X"34",X"06",
		X"DD",X"77",X"05",X"47",X"3A",X"01",X"89",X"FE",X"03",X"DA",X"2D",X"36",X"3A",X"79",X"8D",X"A7",
		X"20",X"32",X"21",X"C7",X"35",X"3A",X"07",X"89",X"E6",X"0F",X"CB",X"3F",X"CD",X"45",X"0C",X"EB",
		X"3A",X"41",X"8D",X"E6",X"07",X"E7",X"4F",X"DD",X"7E",X"06",X"B9",X"CA",X"17",X"36",X"FE",X"14",
		X"D8",X"DD",X"36",X"08",X"01",X"11",X"38",X"38",X"DD",X"CB",X"07",X"4E",X"28",X"03",X"11",X"56",
		X"38",X"C3",X"1E",X"38",X"DD",X"CB",X"07",X"56",X"28",X"08",X"2A",X"6F",X"8D",X"3A",X"7B",X"8D",
		X"18",X"D3",X"DD",X"7E",X"06",X"18",X"D7",X"D7",X"35",X"DF",X"35",X"E7",X"35",X"EF",X"35",X"F7",
		X"35",X"FF",X"35",X"07",X"36",X"0F",X"36",X"09",X"0D",X"11",X"09",X"0D",X"11",X"09",X"0D",X"09",
		X"11",X"0D",X"11",X"0D",X"09",X"0D",X"09",X"11",X"0D",X"09",X"11",X"0D",X"09",X"11",X"0D",X"08",
		X"0B",X"0F",X"12",X"08",X"12",X"0B",X"0F",X"12",X"0F",X"0B",X"08",X"0F",X"12",X"08",X"0B",X"08",
		X"0B",X"0E",X"11",X"0B",X"08",X"11",X"0E",X"11",X"0E",X"0B",X"08",X"0E",X"11",X"0B",X"08",X"08",
		X"0B",X"0F",X"12",X"0A",X"11",X"09",X"0D",X"78",X"FE",X"20",X"D0",X"18",X"40",X"DD",X"CB",X"08",
		X"46",X"C8",X"C3",X"75",X"37",X"DD",X"CB",X"08",X"46",X"C0",X"C3",X"7C",X"35",X"DD",X"7E",X"06",
		X"FE",X"07",X"38",X"E9",X"FE",X"14",X"30",X"ED",X"3A",X"7D",X"8D",X"FE",X"0E",X"38",X"06",X"DD",
		X"7E",X"06",X"FE",X"13",X"D8",X"21",X"6B",X"8D",X"7E",X"A7",X"28",X"02",X"35",X"C9",X"78",X"FE",
		X"80",X"D0",X"EB",X"21",X"8E",X"36",X"3A",X"07",X"89",X"E6",X"07",X"E7",X"12",X"DD",X"CB",X"0B",
		X"46",X"28",X"14",X"21",X"E2",X"8A",X"11",X"18",X"00",X"4A",X"06",X"06",X"7E",X"FE",X"03",X"20",
		X"01",X"0C",X"19",X"10",X"F7",X"0D",X"C0",X"FD",X"21",X"70",X"8B",X"11",X"18",X"00",X"06",X"05",
		X"FD",X"7E",X"00",X"FD",X"B6",X"01",X"0F",X"30",X"0D",X"FD",X"19",X"10",X"F3",X"C9",X"28",X"28",
		X"20",X"20",X"18",X"18",X"10",X"10",X"DD",X"CB",X"07",X"56",X"28",X"13",X"21",X"7B",X"8D",X"34",
		X"21",X"79",X"8D",X"7E",X"A7",X"28",X"08",X"35",X"21",X"75",X"8D",X"77",X"2C",X"36",X"00",X"21",
		X"41",X"8D",X"34",X"20",X"01",X"34",X"4E",X"DD",X"71",X"14",X"21",X"88",X"39",X"DD",X"CB",X"07",
		X"4E",X"28",X"03",X"21",X"94",X"39",X"DD",X"75",X"0C",X"DD",X"74",X"0D",X"DD",X"36",X"0E",X"00",
		X"DD",X"36",X"11",X"28",X"DD",X"36",X"02",X"04",X"CD",X"DE",X"36",X"C3",X"9D",X"37",X"3A",X"07",
		X"89",X"FE",X"10",X"38",X"02",X"3E",X"0E",X"47",X"3A",X"20",X"88",X"87",X"80",X"21",X"37",X"37",
		X"E7",X"DD",X"CB",X"16",X"46",X"28",X"0C",X"3D",X"28",X"16",X"DD",X"CB",X"13",X"46",X"28",X"03",
		X"3D",X"28",X"0D",X"47",X"DD",X"7E",X"06",X"FE",X"09",X"78",X"30",X"04",X"3D",X"28",X"01",X"3D",
		X"47",X"3A",X"01",X"89",X"FE",X"04",X"78",X"30",X"03",X"3E",X"03",X"80",X"21",X"27",X"37",X"E7",
		X"DD",X"B6",X"08",X"DD",X"77",X"08",X"C9",X"00",X"10",X"20",X"30",X"40",X"50",X"60",X"70",X"80",
		X"90",X"A0",X"B0",X"C0",X"D0",X"E0",X"F0",X"01",X"01",X"02",X"02",X"03",X"02",X"04",X"02",X"05",
		X"03",X"05",X"03",X"06",X"03",X"06",X"03",X"07",X"03",X"07",X"03",X"07",X"04",X"07",X"04",X"07",
		X"04",X"07",X"04",X"07",X"04",X"07",X"04",X"DD",X"7E",X"0A",X"ED",X"44",X"47",X"DD",X"7E",X"05",
		X"B8",X"30",X"03",X"DD",X"35",X"06",X"DD",X"86",X"0A",X"DD",X"77",X"05",X"47",X"3A",X"01",X"89",
		X"FE",X"03",X"DA",X"2D",X"36",X"3A",X"0A",X"88",X"FE",X"05",X"28",X"19",X"DD",X"7E",X"06",X"FE",
		X"02",X"D0",X"DD",X"36",X"08",X"00",X"11",X"29",X"38",X"DD",X"CB",X"07",X"4E",X"28",X"03",X"11",
		X"47",X"38",X"C3",X"1E",X"38",X"DD",X"7E",X"06",X"A7",X"C0",X"C3",X"53",X"35",X"FD",X"36",X"00",
		X"01",X"FD",X"36",X"02",X"04",X"FD",X"71",X"14",X"AF",X"FD",X"77",X"07",X"FD",X"77",X"0E",X"DD",
		X"7E",X"05",X"C6",X"80",X"FD",X"77",X"05",X"DD",X"7E",X"03",X"C6",X"80",X"FD",X"77",X"03",X"DD",
		X"7E",X"04",X"D6",X"01",X"FD",X"77",X"04",X"DD",X"7E",X"06",X"C6",X"01",X"FD",X"77",X"06",X"21",
		X"A5",X"38",X"3A",X"20",X"88",X"FE",X"07",X"20",X"03",X"21",X"AD",X"38",X"3A",X"00",X"89",X"FE",
		X"08",X"38",X"02",X"3E",X"07",X"E7",X"3A",X"07",X"89",X"E6",X"01",X"7E",X"28",X"02",X"ED",X"44",
		X"FD",X"77",X"0A",X"DD",X"77",X"0A",X"21",X"B5",X"38",X"DD",X"7E",X"07",X"E6",X"F0",X"0F",X"0F",
		X"0F",X"0F",X"CD",X"45",X"0C",X"DD",X"7E",X"0B",X"A7",X"28",X"03",X"11",X"52",X"39",X"FD",X"77",
		X"0B",X"FD",X"73",X"0C",X"FD",X"72",X"0D",X"FD",X"36",X"11",X"28",X"C3",X"E3",X"0E",X"DD",X"73",
		X"0C",X"DD",X"72",X"0D",X"DD",X"36",X"0E",X"00",X"C9",X"40",X"26",X"07",X"40",X"27",X"07",X"40",
		X"28",X"07",X"40",X"27",X"07",X"FF",X"29",X"38",X"C0",X"26",X"07",X"C0",X"27",X"07",X"C0",X"28",
		X"07",X"C0",X"27",X"07",X"FF",X"38",X"38",X"44",X"26",X"07",X"44",X"27",X"07",X"44",X"28",X"07",
		X"44",X"27",X"07",X"FF",X"47",X"38",X"C4",X"26",X"07",X"C4",X"27",X"07",X"C4",X"28",X"07",X"C4",
		X"27",X"07",X"FF",X"56",X"38",X"CD",X"06",X"40",X"DD",X"35",X"11",X"C0",X"DD",X"34",X"02",X"DD",
		X"CB",X"08",X"86",X"DD",X"E5",X"E1",X"7C",X"FE",X"8B",X"D8",X"7D",X"FE",X"70",X"D8",X"DD",X"35",
		X"04",X"DD",X"35",X"06",X"3A",X"5F",X"8A",X"A7",X"C0",X"21",X"82",X"42",X"0E",X"00",X"59",X"7E",
		X"2B",X"81",X"4F",X"30",X"01",X"1C",X"3E",X"1A",X"BE",X"20",X"F4",X"7B",X"81",X"E6",X"9E",X"C8",
		X"21",X"F0",X"8E",X"34",X"C9",X"10",X"11",X"12",X"13",X"14",X"15",X"16",X"17",X"13",X"14",X"15",
		X"16",X"17",X"17",X"17",X"17",X"CB",X"38",X"DA",X"38",X"E9",X"38",X"F8",X"38",X"07",X"39",X"16",
		X"39",X"25",X"39",X"25",X"39",X"25",X"39",X"34",X"39",X"43",X"39",X"40",X"2D",X"12",X"40",X"02",
		X"0C",X"40",X"3B",X"06",X"40",X"A1",X"E0",X"FF",X"D4",X"38",X"41",X"2D",X"12",X"41",X"02",X"0C",
		X"41",X"3B",X"06",X"41",X"A1",X"E0",X"FF",X"E3",X"38",X"44",X"2D",X"12",X"44",X"02",X"0C",X"44",
		X"3B",X"06",X"44",X"A1",X"E0",X"FF",X"F2",X"38",X"49",X"2D",X"12",X"49",X"02",X"0C",X"49",X"3B",
		X"06",X"49",X"A1",X"E0",X"FF",X"01",X"39",X"4A",X"2D",X"12",X"4A",X"02",X"0C",X"4A",X"3B",X"06",
		X"4A",X"A1",X"E0",X"FF",X"10",X"39",X"41",X"2D",X"12",X"41",X"02",X"0C",X"41",X"3B",X"06",X"41",
		X"A1",X"E0",X"FF",X"1F",X"39",X"44",X"2D",X"12",X"44",X"02",X"0C",X"44",X"3B",X"06",X"44",X"A1",
		X"E0",X"FF",X"2E",X"39",X"4E",X"2D",X"12",X"4E",X"02",X"0C",X"4E",X"3B",X"06",X"4E",X"A1",X"E0",
		X"FF",X"3D",X"39",X"4F",X"2D",X"12",X"4F",X"02",X"0C",X"4F",X"3B",X"06",X"4F",X"A1",X"E0",X"FF",
		X"4C",X"39",X"44",X"2D",X"12",X"44",X"02",X"0C",X"44",X"3B",X"06",X"44",X"A1",X"08",X"4B",X"A1",
		X"08",X"4C",X"A1",X"08",X"4F",X"A1",X"08",X"FF",X"5B",X"39",X"40",X"2A",X"12",X"40",X"2B",X"18",
		X"40",X"29",X"20",X"40",X"1F",X"10",X"FF",X"70",X"39",X"44",X"2A",X"12",X"44",X"2B",X"18",X"44",
		X"29",X"20",X"44",X"1F",X"10",X"FF",X"7F",X"39",X"40",X"26",X"28",X"40",X"29",X"20",X"40",X"1F",
		X"10",X"FF",X"8B",X"39",X"44",X"26",X"28",X"44",X"29",X"20",X"44",X"1F",X"10",X"FF",X"97",X"39",
		X"40",X"2A",X"12",X"40",X"2B",X"18",X"40",X"06",X"10",X"40",X"0B",X"10",X"FF",X"A6",X"39",X"CD",
		X"06",X"40",X"3A",X"07",X"89",X"E6",X"01",X"CA",X"87",X"3B",X"DD",X"7E",X"0A",X"ED",X"44",X"47",
		X"DD",X"7E",X"03",X"B8",X"30",X"03",X"DD",X"35",X"04",X"DD",X"86",X"0A",X"DD",X"77",X"03",X"DD",
		X"46",X"04",X"DD",X"7E",X"07",X"A7",X"28",X"79",X"78",X"FE",X"04",X"38",X"6B",X"FE",X"10",X"D8",
		X"21",X"7D",X"8D",X"7E",X"FE",X"0E",X"30",X"20",X"3A",X"07",X"89",X"FE",X"06",X"30",X"0C",X"3A",
		X"08",X"89",X"FE",X"03",X"38",X"05",X"7E",X"FE",X"08",X"30",X"0D",X"3A",X"20",X"88",X"FE",X"07",
		X"28",X"06",X"DD",X"7E",X"06",X"FE",X"10",X"D0",X"3A",X"75",X"8D",X"A7",X"C0",X"DD",X"7E",X"08",
		X"E6",X"F0",X"C8",X"DD",X"7E",X"15",X"A7",X"28",X"04",X"DD",X"35",X"15",X"C9",X"3A",X"42",X"88",
		X"4F",X"3A",X"1F",X"88",X"47",X"A7",X"79",X"20",X"02",X"ED",X"44",X"0F",X"0F",X"0F",X"E6",X"1F",
		X"4F",X"78",X"A7",X"20",X"02",X"0D",X"0D",X"3A",X"07",X"89",X"47",X"CB",X"47",X"79",X"28",X"02",
		X"C6",X"04",X"DD",X"BE",X"04",X"28",X"25",X"C9",X"DD",X"36",X"02",X"00",X"DD",X"36",X"11",X"20",
		X"C9",X"78",X"FE",X"02",X"D0",X"11",X"D1",X"3B",X"CD",X"1E",X"38",X"DD",X"36",X"02",X"02",X"DD",
		X"36",X"11",X"28",X"C9",X"10",X"15",X"0D",X"1B",X"0F",X"11",X"13",X"1C",X"21",X"42",X"8D",X"34",
		X"FD",X"21",X"E8",X"8B",X"06",X"03",X"11",X"18",X"00",X"FD",X"7E",X"00",X"FD",X"B6",X"01",X"0F",
		X"30",X"05",X"FD",X"19",X"10",X"F3",X"C9",X"DD",X"7E",X"06",X"D6",X"06",X"CB",X"3F",X"E6",X"07",
		X"4F",X"21",X"57",X"3B",X"3A",X"07",X"89",X"CB",X"47",X"28",X"03",X"21",X"47",X"3B",X"79",X"CD",
		X"45",X"0C",X"1A",X"FD",X"77",X"12",X"13",X"1A",X"FD",X"77",X"13",X"FD",X"CB",X"08",X"C6",X"11",
		X"6A",X"39",X"DD",X"CB",X"07",X"4E",X"28",X"03",X"11",X"79",X"39",X"DD",X"7E",X"16",X"E6",X"30",
		X"FE",X"30",X"20",X"03",X"11",X"A0",X"39",X"CD",X"1E",X"38",X"DD",X"7E",X"08",X"D6",X"10",X"DD",
		X"77",X"08",X"FD",X"36",X"00",X"01",X"FD",X"36",X"02",X"0B",X"FD",X"36",X"07",X"01",X"3A",X"50",
		X"8F",X"A7",X"11",X"DD",X"3B",X"28",X"0D",X"11",X"3B",X"43",X"3A",X"07",X"89",X"CB",X"57",X"28",
		X"03",X"11",X"41",X"43",X"FD",X"73",X"0C",X"FD",X"72",X"0D",X"FD",X"36",X"0E",X"00",X"FD",X"36",
		X"16",X"00",X"FD",X"36",X"11",X"13",X"DD",X"E5",X"E1",X"FD",X"75",X"14",X"FD",X"74",X"15",X"21",
		X"6C",X"8D",X"34",X"7E",X"E6",X"07",X"57",X"21",X"37",X"3B",X"3A",X"07",X"89",X"CB",X"47",X"28",
		X"03",X"21",X"3F",X"3B",X"7A",X"E7",X"DD",X"77",X"15",X"C9",X"00",X"01",X"01",X"04",X"04",X"04",
		X"07",X"0A",X"0D",X"0D",X"0D",X"0D",X"0D",X"20",X"1C",X"18",X"20",X"28",X"30",X"18",X"30",X"20",
		X"22",X"24",X"26",X"28",X"30",X"28",X"30",X"67",X"3B",X"69",X"3B",X"6B",X"3B",X"6D",X"3B",X"6F",
		X"3B",X"71",X"3B",X"73",X"3B",X"75",X"3B",X"77",X"3B",X"79",X"3B",X"7B",X"3B",X"7D",X"3B",X"7F",
		X"3B",X"81",X"3B",X"83",X"3B",X"85",X"3B",X"40",X"48",X"40",X"48",X"40",X"40",X"40",X"44",X"40",
		X"48",X"40",X"50",X"40",X"58",X"40",X"30",X"40",X"20",X"40",X"20",X"40",X"1C",X"40",X"1C",X"40",
		X"1C",X"40",X"18",X"40",X"18",X"40",X"38",X"DD",X"CB",X"08",X"46",X"C2",X"BA",X"39",X"DD",X"7E",
		X"03",X"DD",X"86",X"0A",X"30",X"03",X"DD",X"34",X"04",X"DD",X"77",X"03",X"DD",X"46",X"04",X"DD",
		X"7E",X"07",X"A7",X"CA",X"CA",X"3B",X"78",X"FE",X"1D",X"30",X"03",X"C3",X"E0",X"39",X"DD",X"34",
		X"02",X"AF",X"DD",X"77",X"00",X"DD",X"36",X"01",X"01",X"DD",X"CB",X"08",X"86",X"DD",X"36",X"09",
		X"20",X"DD",X"77",X"14",X"11",X"29",X"38",X"C3",X"1E",X"38",X"78",X"FE",X"1B",X"D4",X"53",X"35",
		X"C9",X"40",X"34",X"07",X"40",X"33",X"08",X"40",X"32",X"09",X"40",X"31",X"20",X"40",X"00",X"F0",
		X"FF",X"DD",X"3B",X"CD",X"06",X"40",X"DD",X"CB",X"08",X"46",X"20",X"24",X"DD",X"7E",X"05",X"DD",
		X"86",X"09",X"30",X"03",X"DD",X"34",X"06",X"DD",X"77",X"05",X"47",X"DD",X"7E",X"06",X"FE",X"1F",
		X"D8",X"18",X"38",X"DD",X"34",X"02",X"DD",X"36",X"11",X"20",X"3E",X"28",X"32",X"5E",X"8D",X"C9",
		X"DD",X"7E",X"0A",X"ED",X"44",X"47",X"DD",X"7E",X"05",X"B8",X"30",X"03",X"DD",X"35",X"06",X"DD",
		X"86",X"0A",X"DD",X"77",X"05",X"47",X"DD",X"6E",X"14",X"DD",X"66",X"15",X"E5",X"FD",X"E1",X"FD",
		X"77",X"05",X"DD",X"7E",X"06",X"FD",X"77",X"06",X"E6",X"1F",X"C0",X"21",X"03",X"89",X"34",X"21",
		X"40",X"8D",X"35",X"2E",X"7D",X"34",X"DD",X"7E",X"07",X"E6",X"F0",X"CA",X"53",X"35",X"CD",X"53",
		X"35",X"3A",X"7E",X"8D",X"A7",X"C0",X"21",X"76",X"8D",X"34",X"7E",X"FE",X"02",X"D8",X"2D",X"AF",
		X"77",X"32",X"20",X"8F",X"32",X"6D",X"8D",X"32",X"6E",X"8D",X"3E",X"02",X"32",X"07",X"8D",X"32",
		X"7E",X"8D",X"3A",X"1F",X"88",X"A7",X"C0",X"3A",X"01",X"89",X"FE",X"10",X"D0",X"11",X"D5",X"01",
		X"01",X"12",X"00",X"1A",X"1B",X"80",X"47",X"0D",X"20",X"F9",X"FE",X"55",X"C8",X"21",X"ED",X"89",
		X"34",X"C9",X"CD",X"06",X"40",X"DD",X"35",X"11",X"C0",X"FD",X"21",X"30",X"8C",X"11",X"18",X"00",
		X"06",X"04",X"CD",X"AE",X"3C",X"FD",X"19",X"10",X"F9",X"DD",X"36",X"11",X"10",X"C9",X"FD",X"7E",
		X"00",X"FD",X"B6",X"01",X"0F",X"C0",X"FD",X"36",X"01",X"01",X"AF",X"FD",X"36",X"02",X"10",X"21",
		X"0F",X"3D",X"FD",X"75",X"0C",X"FD",X"74",X"0D",X"FD",X"77",X"0E",X"DD",X"36",X"02",X"06",X"DD",
		X"36",X"08",X"01",X"DD",X"36",X"0A",X"E8",X"11",X"38",X"38",X"CD",X"1E",X"38",X"DD",X"7E",X"04",
		X"D6",X"01",X"FD",X"77",X"04",X"DD",X"7E",X"03",X"FD",X"77",X"03",X"DD",X"7E",X"06",X"C6",X"01",
		X"FD",X"77",X"06",X"DD",X"7E",X"05",X"FD",X"77",X"05",X"FD",X"36",X"08",X"01",X"FD",X"36",X"0A",
		X"E8",X"CD",X"3C",X"40",X"FD",X"E5",X"E1",X"DD",X"75",X"14",X"DD",X"74",X"15",X"F1",X"C9",X"40",
		X"83",X"10",X"40",X"89",X"10",X"FF",X"0F",X"3D",X"06",X"20",X"DD",X"4E",X"17",X"3A",X"45",X"8D",
		X"A7",X"28",X"18",X"DD",X"4E",X"12",X"0C",X"28",X"12",X"FE",X"04",X"38",X"02",X"3E",X"03",X"47",
		X"C6",X"06",X"4F",X"11",X"0F",X"03",X"83",X"5F",X"FF",X"06",X"38",X"DD",X"70",X"11",X"79",X"DD",
		X"CB",X"07",X"4E",X"28",X"0B",X"0C",X"3A",X"45",X"8D",X"A7",X"79",X"28",X"03",X"3E",X"03",X"81",
		X"21",X"D3",X"3D",X"CD",X"45",X"0C",X"CD",X"1E",X"38",X"DD",X"34",X"02",X"CD",X"06",X"40",X"DD",
		X"35",X"11",X"C0",X"DD",X"7E",X"16",X"FE",X"07",X"CA",X"99",X"3D",X"4F",X"A7",X"28",X"01",X"3D",
		X"11",X"12",X"03",X"83",X"5F",X"FF",X"21",X"49",X"3E",X"79",X"FE",X"04",X"20",X"0A",X"CD",X"45",
		X"0C",X"CD",X"1E",X"38",X"DD",X"36",X"11",X"30",X"0C",X"DD",X"71",X"13",X"DD",X"34",X"02",X"CD",
		X"06",X"40",X"DD",X"35",X"11",X"C0",X"C3",X"53",X"35",X"21",X"76",X"40",X"DD",X"7E",X"07",X"E6",
		X"03",X"3D",X"CD",X"45",X"0C",X"CD",X"1E",X"38",X"DD",X"36",X"09",X"40",X"DD",X"36",X"02",X"0F",
		X"C3",X"D6",X"0E",X"BB",X"3D",X"C1",X"3D",X"C7",X"3D",X"CD",X"3D",X"42",X"30",X"F0",X"FF",X"BB",
		X"3D",X"41",X"30",X"F0",X"FF",X"C1",X"3D",X"49",X"30",X"F0",X"FF",X"C7",X"3D",X"40",X"30",X"F0",
		X"FF",X"CD",X"3D",X"EF",X"3D",X"EF",X"3D",X"EF",X"3D",X"FB",X"3D",X"07",X"3E",X"7A",X"40",X"8F",
		X"40",X"13",X"3E",X"1C",X"3E",X"25",X"3E",X"25",X"3E",X"2E",X"3E",X"37",X"3E",X"40",X"3E",X"44",
		X"34",X"05",X"44",X"33",X"06",X"44",X"32",X"07",X"44",X"31",X"12",X"40",X"34",X"05",X"40",X"33",
		X"06",X"40",X"32",X"07",X"40",X"31",X"12",X"40",X"34",X"05",X"40",X"33",X"06",X"40",X"32",X"07",
		X"40",X"31",X"12",X"80",X"01",X"05",X"40",X"1D",X"05",X"43",X"39",X"28",X"80",X"01",X"04",X"40",
		X"1D",X"04",X"42",X"39",X"28",X"80",X"01",X"03",X"40",X"1D",X"03",X"4F",X"3A",X"38",X"84",X"01",
		X"05",X"44",X"1D",X"05",X"43",X"39",X"28",X"84",X"01",X"04",X"44",X"1D",X"04",X"42",X"39",X"28",
		X"84",X"01",X"03",X"44",X"1D",X"03",X"4F",X"3A",X"38",X"5D",X"3E",X"5D",X"3E",X"5D",X"3E",X"5D",
		X"3E",X"5D",X"3E",X"63",X"3E",X"66",X"3E",X"66",X"3E",X"66",X"3E",X"66",X"3E",X"42",X"37",X"40",
		X"43",X"39",X"40",X"42",X"39",X"40",X"4F",X"3B",X"48",X"DD",X"35",X"11",X"C0",X"DD",X"6E",X"14",
		X"DD",X"66",X"15",X"2C",X"2C",X"7E",X"FE",X"05",X"DA",X"53",X"35",X"FE",X"07",X"D2",X"53",X"35",
		X"2C",X"7E",X"DD",X"77",X"03",X"2C",X"7E",X"3D",X"DD",X"77",X"04",X"2C",X"7E",X"DD",X"77",X"05",
		X"2C",X"7E",X"DD",X"77",X"06",X"DD",X"36",X"15",X"00",X"DD",X"34",X"02",X"CD",X"06",X"40",X"DD",
		X"CB",X"01",X"46",X"C2",X"1D",X"3F",X"DD",X"6E",X"12",X"DD",X"66",X"13",X"DD",X"7E",X"05",X"85",
		X"DD",X"77",X"05",X"30",X"03",X"DD",X"34",X"06",X"DD",X"CB",X"08",X"46",X"28",X"43",X"7C",X"D6",
		X"02",X"38",X"35",X"67",X"DD",X"7E",X"03",X"94",X"DD",X"77",X"03",X"30",X"03",X"DD",X"35",X"04",
		X"DD",X"74",X"13",X"DD",X"7E",X"06",X"E6",X"1F",X"FE",X"1A",X"D8",X"DD",X"7E",X"05",X"FE",X"A0",
		X"D0",X"11",X"B4",X"40",X"CD",X"1E",X"38",X"DD",X"36",X"11",X"0A",X"DD",X"36",X"02",X"02",X"DD",
		X"36",X"00",X"00",X"DD",X"36",X"01",X"01",X"C9",X"DD",X"CB",X"08",X"86",X"AF",X"DD",X"77",X"13",
		X"C9",X"DD",X"34",X"16",X"DD",X"7E",X"16",X"E6",X"03",X"C8",X"7C",X"C6",X"01",X"DD",X"77",X"13",
		X"DD",X"86",X"03",X"DD",X"77",X"03",X"30",X"03",X"DD",X"34",X"04",X"18",X"B6",X"DD",X"6E",X"12",
		X"DD",X"66",X"13",X"7E",X"4F",X"FE",X"EE",X"20",X"01",X"23",X"46",X"DD",X"7E",X"05",X"90",X"DD",
		X"77",X"05",X"30",X"03",X"DD",X"35",X"06",X"23",X"7E",X"DD",X"86",X"03",X"DD",X"77",X"03",X"30",
		X"03",X"DD",X"34",X"04",X"23",X"79",X"FE",X"EE",X"20",X"03",X"2B",X"2B",X"2B",X"DD",X"75",X"12",
		X"DD",X"74",X"13",X"DD",X"7E",X"04",X"FE",X"1E",X"D8",X"C3",X"E1",X"3E",X"21",X"72",X"40",X"DD",
		X"7E",X"07",X"E6",X"03",X"3D",X"CD",X"45",X"0C",X"CD",X"1E",X"38",X"DD",X"36",X"09",X"40",X"DD",
		X"34",X"02",X"CD",X"06",X"40",X"DD",X"35",X"11",X"C0",X"DD",X"34",X"02",X"CD",X"06",X"40",X"CD",
		X"D5",X"3F",X"D8",X"21",X"A4",X"40",X"DD",X"7E",X"07",X"E6",X"03",X"3D",X"CD",X"45",X"0C",X"CD",
		X"1E",X"38",X"DD",X"36",X"02",X"02",X"DD",X"36",X"11",X"20",X"CD",X"DA",X"0E",X"21",X"40",X"8D",
		X"35",X"21",X"01",X"89",X"DD",X"CB",X"0B",X"46",X"20",X"07",X"7E",X"A7",X"C8",X"35",X"C3",X"C9",
		X"34",X"36",X"00",X"3E",X"01",X"CD",X"C9",X"34",X"01",X"8B",X"42",X"2E",X"00",X"65",X"0A",X"FE",
		X"C8",X"28",X"08",X"84",X"30",X"01",X"2C",X"67",X"0B",X"18",X"F3",X"95",X"FE",X"C0",X"C8",X"3E",
		X"01",X"32",X"EB",X"89",X"C9",X"DD",X"7E",X"03",X"DD",X"86",X"09",X"30",X"03",X"DD",X"34",X"04",
		X"DD",X"77",X"03",X"DD",X"7E",X"04",X"FE",X"1E",X"C9",X"11",X"80",X"77",X"01",X"10",X"00",X"1A",
		X"1B",X"80",X"47",X"0D",X"20",X"F9",X"CB",X"40",X"20",X"07",X"CB",X"68",X"28",X"03",X"CB",X"78",
		X"C0",X"21",X"39",X"8A",X"34",X"C9",X"DD",X"7E",X"0E",X"A7",X"28",X"04",X"DD",X"35",X"0E",X"C9",
		X"DD",X"6E",X"0C",X"DD",X"66",X"0D",X"7E",X"FE",X"FF",X"28",X"15",X"DD",X"77",X"10",X"23",X"7E",
		X"DD",X"77",X"0F",X"23",X"7E",X"DD",X"77",X"0E",X"23",X"DD",X"75",X"0C",X"DD",X"74",X"0D",X"C9",
		X"23",X"7E",X"DD",X"77",X"0C",X"23",X"7E",X"DD",X"77",X"0D",X"18",X"D4",X"FD",X"7E",X"0E",X"A7",
		X"28",X"04",X"FD",X"35",X"0E",X"C9",X"FD",X"6E",X"0C",X"FD",X"66",X"0D",X"7E",X"FE",X"FF",X"28",
		X"15",X"FD",X"77",X"10",X"23",X"7E",X"FD",X"77",X"0F",X"23",X"7E",X"FD",X"77",X"0E",X"23",X"FD",
		X"75",X"0C",X"FD",X"74",X"0D",X"C9",X"23",X"7E",X"FD",X"77",X"0C",X"23",X"7E",X"FD",X"77",X"0D",
		X"18",X"D4",X"7A",X"40",X"8F",X"40",X"86",X"40",X"9B",X"40",X"80",X"01",X"08",X"40",X"1D",X"08",
		X"80",X"01",X"08",X"40",X"1D",X"08",X"40",X"01",X"08",X"80",X"1D",X"08",X"FF",X"86",X"40",X"84",
		X"01",X"08",X"44",X"1D",X"08",X"84",X"01",X"08",X"44",X"1D",X"08",X"44",X"01",X"08",X"84",X"1D",
		X"08",X"FF",X"9B",X"40",X"A8",X"40",X"AE",X"40",X"40",X"19",X"28",X"40",X"19",X"38",X"44",X"19",
		X"28",X"44",X"19",X"30",X"45",X"34",X"05",X"45",X"33",X"05",X"FF",X"B4",X"40",X"DD",X"21",X"30",
		X"8C",X"11",X"18",X"00",X"06",X"04",X"D9",X"CD",X"D0",X"40",X"D9",X"DD",X"19",X"10",X"F7",X"C9",
		X"DD",X"7E",X"00",X"DD",X"B6",X"01",X"0F",X"D0",X"DD",X"7E",X"02",X"E6",X"1F",X"FE",X"11",X"D0",
		X"EF",X"03",X"41",X"37",X"41",X"6F",X"41",X"79",X"41",X"79",X"41",X"79",X"41",X"79",X"41",X"79",
		X"41",X"7A",X"41",X"8D",X"41",X"79",X"41",X"21",X"42",X"50",X"43",X"64",X"43",X"78",X"43",X"78",
		X"43",X"78",X"43",X"CD",X"06",X"40",X"DD",X"35",X"11",X"C0",X"DD",X"34",X"02",X"DD",X"36",X"13",
		X"00",X"3A",X"5F",X"8A",X"A7",X"C0",X"21",X"7F",X"55",X"06",X"38",X"AF",X"57",X"5A",X"7E",X"E6",
		X"0F",X"83",X"5F",X"30",X"01",X"14",X"23",X"10",X"F5",X"3E",X"67",X"BB",X"20",X"04",X"3E",X"01",
		X"92",X"C8",X"21",X"38",X"8A",X"34",X"C9",X"CD",X"06",X"40",X"DD",X"7E",X"0A",X"ED",X"44",X"47",
		X"DD",X"7E",X"03",X"B8",X"30",X"03",X"DD",X"35",X"04",X"DD",X"86",X"0A",X"DD",X"77",X"03",X"47",
		X"DD",X"7E",X"04",X"FE",X"03",X"D0",X"DD",X"7E",X"17",X"3C",X"32",X"1D",X"8D",X"3D",X"DD",X"36",
		X"02",X"02",X"DD",X"36",X"11",X"18",X"21",X"B1",X"41",X"CD",X"45",X"0C",X"C3",X"1E",X"38",X"CD",
		X"06",X"40",X"DD",X"35",X"11",X"C0",X"C3",X"53",X"35",X"C9",X"DD",X"7E",X"17",X"21",X"B1",X"41",
		X"CD",X"45",X"0C",X"CD",X"1E",X"38",X"DD",X"36",X"11",X"30",X"DD",X"34",X"02",X"CD",X"06",X"40",
		X"DD",X"35",X"11",X"C0",X"DD",X"7E",X"16",X"4F",X"A7",X"28",X"01",X"3D",X"11",X"12",X"03",X"83",
		X"5F",X"FF",X"DD",X"36",X"11",X"01",X"0C",X"DD",X"71",X"13",X"DD",X"36",X"02",X"02",X"C3",X"6F",
		X"41",X"BB",X"41",X"CA",X"41",X"D9",X"41",X"E8",X"41",X"F7",X"41",X"44",X"34",X"05",X"44",X"33",
		X"06",X"44",X"32",X"07",X"44",X"31",X"08",X"43",X"37",X"38",X"41",X"34",X"05",X"41",X"33",X"06",
		X"41",X"32",X"07",X"41",X"31",X"08",X"43",X"37",X"38",X"49",X"34",X"05",X"49",X"33",X"06",X"49",
		X"32",X"07",X"49",X"31",X"08",X"43",X"37",X"38",X"40",X"34",X"05",X"40",X"33",X"06",X"40",X"32",
		X"07",X"40",X"31",X"08",X"48",X"37",X"38",X"47",X"34",X"05",X"47",X"33",X"06",X"47",X"32",X"07",
		X"47",X"31",X"12",X"44",X"26",X"09",X"44",X"27",X"09",X"44",X"28",X"09",X"44",X"27",X"09",X"FF",
		X"03",X"42",X"C4",X"26",X"09",X"C4",X"27",X"09",X"C4",X"28",X"09",X"C4",X"27",X"09",X"FF",X"12",
		X"42",X"CD",X"06",X"40",X"DD",X"CB",X"08",X"46",X"20",X"1A",X"CD",X"3E",X"34",X"DD",X"7E",X"06",
		X"E6",X"1F",X"FE",X"14",X"38",X"5A",X"DD",X"36",X"08",X"01",X"11",X"12",X"42",X"AF",X"32",X"4B",
		X"8D",X"C3",X"1E",X"38",X"CD",X"F2",X"34",X"DD",X"7E",X"06",X"E6",X"1F",X"FE",X"0A",X"30",X"40",
		X"47",X"3A",X"01",X"89",X"FE",X"02",X"38",X"0E",X"DD",X"36",X"08",X"00",X"11",X"03",X"42",X"3E",
		X"FF",X"32",X"4B",X"8D",X"18",X"DB",X"78",X"FE",X"02",X"D0",X"CD",X"53",X"35",X"11",X"B9",X"0B",
		X"21",X"83",X"42",X"1A",X"86",X"20",X"07",X"1B",X"23",X"7E",X"3C",X"C8",X"18",X"F5",X"21",X"3A",
		X"8A",X"34",X"C9",X"E0",X"59",X"78",X"FA",X"C6",X"7A",X"B5",X"7A",X"B2",X"7A",X"AD",X"7A",X"FF",
		X"FE",X"05",X"D8",X"21",X"5B",X"8D",X"7E",X"A7",X"20",X"2F",X"2B",X"7E",X"A7",X"28",X"02",X"35",
		X"C9",X"3A",X"01",X"89",X"FE",X"08",X"11",X"18",X"00",X"38",X"15",X"FD",X"21",X"E0",X"8A",X"3A",
		X"5C",X"8D",X"47",X"4F",X"FD",X"7E",X"04",X"FE",X"07",X"28",X"05",X"FD",X"19",X"10",X"F5",X"C9",
		X"3A",X"5D",X"8D",X"32",X"5A",X"8D",X"32",X"5B",X"8D",X"FD",X"21",X"48",X"8C",X"06",X"03",X"CD",
		X"DA",X"42",X"11",X"18",X"00",X"FD",X"19",X"10",X"F6",X"C9",X"FD",X"7E",X"00",X"FD",X"B6",X"01",
		X"0F",X"D8",X"FD",X"36",X"00",X"01",X"FD",X"36",X"02",X"0D",X"DD",X"E5",X"E1",X"FD",X"E5",X"D1",
		X"2C",X"2C",X"2C",X"1C",X"1C",X"1C",X"01",X"04",X"00",X"ED",X"B0",X"3E",X"2A",X"FD",X"77",X"09",
		X"ED",X"44",X"FD",X"77",X"0A",X"21",X"2D",X"43",X"3A",X"07",X"89",X"CB",X"3F",X"3D",X"E6",X"03",
		X"CD",X"45",X"0C",X"CD",X"75",X"5C",X"AF",X"32",X"5B",X"8D",X"11",X"47",X"43",X"CD",X"1E",X"38",
		X"DD",X"36",X"11",X"30",X"FD",X"36",X"11",X"04",X"DD",X"34",X"02",X"F1",X"C9",X"35",X"43",X"41",
		X"43",X"3B",X"43",X"41",X"43",X"46",X"1C",X"F0",X"FF",X"35",X"43",X"46",X"1C",X"F0",X"FF",X"3B",
		X"43",X"47",X"1C",X"F0",X"FF",X"41",X"43",X"44",X"2C",X"30",X"44",X"20",X"F0",X"FF",X"4A",X"43",
		X"CD",X"06",X"40",X"DD",X"35",X"11",X"C0",X"DD",X"35",X"02",X"DD",X"CB",X"08",X"46",X"CA",X"5C",
		X"42",X"C3",X"3A",X"42",X"DD",X"7E",X"11",X"A7",X"28",X"04",X"DD",X"35",X"11",X"C9",X"CD",X"06",
		X"40",X"CD",X"D5",X"3F",X"D8",X"C3",X"53",X"35",X"C9",X"10",X"11",X"12",X"13",X"14",X"15",X"16",
		X"17",X"06",X"1D",X"3A",X"20",X"89",X"2A",X"43",X"8F",X"ED",X"5B",X"45",X"8F",X"A7",X"28",X"07",
		X"2A",X"B8",X"88",X"ED",X"5B",X"BA",X"88",X"1A",X"FE",X"10",X"28",X"22",X"FE",X"FF",X"28",X"2E",
		X"77",X"13",X"23",X"10",X"F2",X"23",X"23",X"23",X"3A",X"20",X"89",X"A7",X"20",X"08",X"22",X"43",
		X"8F",X"ED",X"53",X"45",X"8F",X"C9",X"22",X"B8",X"88",X"ED",X"53",X"BA",X"88",X"C9",X"13",X"1A",
		X"4F",X"85",X"30",X"01",X"24",X"6F",X"13",X"78",X"91",X"47",X"20",X"CB",X"18",X"D7",X"13",X"1A",
		X"6F",X"13",X"1A",X"67",X"13",X"1A",X"4F",X"3A",X"B7",X"88",X"81",X"32",X"B7",X"88",X"13",X"18",
		X"C7",X"10",X"10",X"63",X"31",X"4F",X"4F",X"3C",X"75",X"10",X"07",X"10",X"0F",X"46",X"C6",X"30",
		X"3D",X"81",X"3C",X"75",X"10",X"07",X"10",X"10",X"2E",X"32",X"42",X"BD",X"3C",X"75",X"10",X"07",
		X"10",X"0F",X"46",X"2E",X"32",X"3D",X"81",X"3C",X"75",X"10",X"07",X"10",X"10",X"33",X"30",X"42",
		X"BD",X"3C",X"75",X"10",X"07",X"10",X"11",X"6D",X"58",X"58",X"3C",X"75",X"10",X"07",X"10",X"13",
		X"71",X"3C",X"75",X"10",X"07",X"10",X"13",X"71",X"3C",X"75",X"10",X"07",X"10",X"14",X"3C",X"75",
		X"10",X"07",X"10",X"14",X"3C",X"75",X"10",X"07",X"10",X"14",X"3C",X"75",X"10",X"07",X"10",X"14",
		X"3C",X"75",X"10",X"07",X"10",X"14",X"3C",X"75",X"10",X"07",X"10",X"14",X"3C",X"75",X"10",X"07",
		X"10",X"14",X"3C",X"75",X"10",X"07",X"10",X"14",X"3C",X"75",X"10",X"07",X"10",X"14",X"3C",X"75",
		X"10",X"07",X"10",X"14",X"3C",X"75",X"10",X"07",X"10",X"14",X"3C",X"75",X"10",X"07",X"10",X"13",
		X"71",X"3C",X"75",X"10",X"07",X"10",X"14",X"3C",X"75",X"10",X"07",X"10",X"14",X"3C",X"75",X"10",
		X"07",X"10",X"13",X"71",X"3C",X"75",X"10",X"07",X"10",X"14",X"3C",X"75",X"10",X"07",X"10",X"14",
		X"3C",X"75",X"10",X"07",X"10",X"13",X"71",X"3C",X"75",X"10",X"07",X"10",X"13",X"71",X"3C",X"75",
		X"10",X"07",X"10",X"13",X"71",X"3C",X"75",X"10",X"07",X"10",X"07",X"57",X"67",X"4C",X"55",X"67",
		X"72",X"55",X"67",X"4C",X"4C",X"31",X"4F",X"4F",X"3C",X"75",X"10",X"07",X"10",X"06",X"71",X"57",
		X"6B",X"73",X"68",X"6B",X"73",X"68",X"6B",X"73",X"C6",X"30",X"3D",X"81",X"3C",X"75",X"10",X"07",
		X"10",X"07",X"57",X"6A",X"39",X"67",X"6A",X"39",X"67",X"6A",X"39",X"2E",X"32",X"42",X"BD",X"3C",
		X"75",X"10",X"07",X"10",X"07",X"66",X"69",X"3A",X"66",X"69",X"3A",X"66",X"69",X"3A",X"2E",X"32",
		X"3D",X"81",X"3C",X"75",X"10",X"07",X"10",X"10",X"33",X"30",X"42",X"BD",X"3C",X"75",X"10",X"07",
		X"10",X"11",X"6D",X"58",X"58",X"3C",X"75",X"10",X"07",X"10",X"14",X"3C",X"75",X"10",X"07",X"10",
		X"13",X"71",X"3C",X"75",X"10",X"07",X"10",X"01",X"A5",X"A4",X"10",X"11",X"3C",X"75",X"10",X"07",
		X"10",X"01",X"A4",X"A5",X"10",X"11",X"3C",X"75",X"10",X"07",X"10",X"01",X"0C",X"3B",X"10",X"10",
		X"71",X"3C",X"75",X"10",X"07",X"10",X"01",X"0C",X"3B",X"10",X"11",X"3C",X"75",X"10",X"07",X"10",
		X"01",X"0E",X"0F",X"10",X"11",X"3C",X"75",X"10",X"07",X"10",X"01",X"0E",X"0F",X"10",X"04",X"87",
		X"87",X"10",X"0B",X"3C",X"75",X"10",X"07",X"10",X"01",X"0C",X"0C",X"10",X"04",X"9B",X"9D",X"88",
		X"10",X"0A",X"3C",X"75",X"10",X"07",X"10",X"01",X"0C",X"0C",X"10",X"04",X"9C",X"82",X"88",X"10",
		X"0A",X"3C",X"75",X"10",X"07",X"10",X"01",X"0C",X"0C",X"10",X"04",X"79",X"79",X"88",X"10",X"0A",
		X"3C",X"75",X"10",X"07",X"10",X"01",X"0C",X"0C",X"10",X"04",X"9C",X"82",X"87",X"10",X"0A",X"3C",
		X"75",X"10",X"07",X"10",X"01",X"0C",X"0C",X"10",X"04",X"85",X"76",X"87",X"10",X"0A",X"3C",X"75",
		X"10",X"07",X"10",X"01",X"0C",X"0D",X"10",X"04",X"9C",X"79",X"87",X"10",X"0A",X"3C",X"75",X"10",
		X"07",X"10",X"07",X"9C",X"76",X"9B",X"10",X"0A",X"3C",X"75",X"10",X"07",X"10",X"07",X"85",X"76",
		X"9B",X"10",X"0A",X"3C",X"75",X"10",X"07",X"10",X"07",X"85",X"76",X"9D",X"88",X"10",X"09",X"3C",
		X"75",X"10",X"07",X"10",X"07",X"7E",X"7B",X"8F",X"8C",X"10",X"08",X"8B",X"3C",X"75",X"10",X"07",
		X"10",X"07",X"7F",X"7B",X"7C",X"76",X"87",X"10",X"02",X"89",X"86",X"10",X"02",X"86",X"8A",X"3C",
		X"75",X"10",X"07",X"10",X"07",X"85",X"7E",X"7B",X"7C",X"76",X"91",X"83",X"84",X"9E",X"92",X"96",
		X"9E",X"38",X"3C",X"75",X"10",X"07",X"10",X"07",X"9C",X"8E",X"7A",X"78",X"76",X"93",X"9F",X"94",
		X"97",X"94",X"99",X"97",X"97",X"3C",X"75",X"10",X"07",X"10",X"07",X"7E",X"7A",X"7A",X"8E",X"76",
		X"93",X"64",X"98",X"98",X"95",X"95",X"98",X"95",X"3C",X"75",X"10",X"07",X"10",X"14",X"3C",X"75",
		X"10",X"07",X"10",X"14",X"3C",X"75",X"10",X"07",X"10",X"14",X"3C",X"75",X"10",X"07",X"10",X"14",
		X"3C",X"75",X"10",X"07",X"10",X"14",X"3C",X"75",X"10",X"07",X"10",X"14",X"3C",X"75",X"10",X"07",
		X"10",X"14",X"3C",X"75",X"10",X"07",X"10",X"14",X"3C",X"75",X"10",X"07",X"10",X"13",X"71",X"3C",
		X"75",X"10",X"07",X"10",X"14",X"3C",X"75",X"10",X"07",X"10",X"14",X"3C",X"75",X"10",X"07",X"10",
		X"14",X"3C",X"75",X"10",X"07",X"10",X"13",X"71",X"3C",X"75",X"10",X"07",X"10",X"14",X"3C",X"75",
		X"10",X"07",X"10",X"14",X"3C",X"75",X"10",X"07",X"10",X"14",X"3C",X"75",X"10",X"07",X"10",X"14",
		X"3C",X"75",X"10",X"07",X"10",X"14",X"3C",X"75",X"10",X"07",X"10",X"14",X"3C",X"75",X"10",X"07",
		X"10",X"14",X"3C",X"75",X"10",X"07",X"10",X"14",X"3C",X"75",X"10",X"07",X"10",X"14",X"3C",X"75",
		X"10",X"07",X"10",X"14",X"3C",X"75",X"10",X"07",X"10",X"14",X"3C",X"75",X"10",X"07",X"10",X"14",
		X"3C",X"75",X"10",X"07",X"10",X"14",X"3C",X"75",X"10",X"07",X"10",X"14",X"3C",X"75",X"10",X"07",
		X"10",X"14",X"3C",X"75",X"10",X"07",X"10",X"03",X"E6",X"E7",X"57",X"72",X"67",X"72",X"4C",X"55",
		X"55",X"67",X"72",X"4C",X"55",X"67",X"72",X"4C",X"55",X"67",X"72",X"4C",X"63",X"31",X"4F",X"4F",
		X"3C",X"75",X"10",X"03",X"E4",X"E5",X"57",X"72",X"6B",X"73",X"73",X"68",X"68",X"6B",X"73",X"73",
		X"68",X"6B",X"73",X"73",X"68",X"6B",X"73",X"73",X"2E",X"30",X"3D",X"81",X"3C",X"75",X"10",X"03",
		X"E6",X"E7",X"57",X"67",X"6A",X"39",X"39",X"67",X"67",X"6A",X"39",X"39",X"67",X"6A",X"39",X"39",
		X"67",X"6A",X"39",X"39",X"2E",X"32",X"42",X"BD",X"3C",X"75",X"10",X"03",X"A8",X"A9",X"A2",X"A1",
		X"69",X"3A",X"3A",X"66",X"65",X"69",X"3A",X"3A",X"66",X"69",X"3A",X"3A",X"66",X"69",X"3A",X"3A",
		X"2E",X"32",X"3D",X"81",X"3C",X"75",X"10",X"03",X"AA",X"AB",X"10",X"12",X"33",X"30",X"42",X"BD",
		X"3C",X"75",X"10",X"03",X"AF",X"37",X"37",X"37",X"34",X"10",X"10",X"6D",X"58",X"58",X"3C",X"75",
		X"10",X"03",X"87",X"87",X"10",X"16",X"3C",X"75",X"10",X"03",X"9B",X"9D",X"88",X"10",X"15",X"3C",
		X"75",X"10",X"03",X"9C",X"82",X"88",X"10",X"15",X"3C",X"75",X"10",X"03",X"79",X"79",X"88",X"10",
		X"15",X"3C",X"75",X"10",X"03",X"9C",X"82",X"87",X"10",X"14",X"71",X"3C",X"75",X"10",X"03",X"85",
		X"76",X"87",X"10",X"15",X"3C",X"75",X"10",X"03",X"9C",X"76",X"87",X"10",X"15",X"3C",X"75",X"10",
		X"03",X"9C",X"79",X"9B",X"10",X"15",X"3C",X"75",X"10",X"03",X"79",X"76",X"87",X"10",X"14",X"71",
		X"3C",X"75",X"10",X"03",X"80",X"8D",X"10",X"16",X"3C",X"75",X"10",X"03",X"80",X"76",X"87",X"10",
		X"15",X"3C",X"75",X"10",X"03",X"85",X"76",X"9B",X"10",X"15",X"3C",X"75",X"10",X"03",X"85",X"82",
		X"9B",X"10",X"15",X"3C",X"75",X"10",X"03",X"9C",X"79",X"9B",X"10",X"15",X"3C",X"75",X"10",X"03",
		X"9C",X"79",X"9D",X"88",X"10",X"14",X"3C",X"75",X"10",X"03",X"85",X"76",X"76",X"87",X"10",X"14",
		X"3C",X"75",X"10",X"03",X"7E",X"7B",X"90",X"8F",X"8C",X"10",X"13",X"3C",X"75",X"10",X"03",X"7F",
		X"7B",X"7C",X"76",X"76",X"87",X"10",X"11",X"8B",X"3C",X"75",X"10",X"03",X"85",X"79",X"76",X"76",
		X"79",X"9D",X"88",X"10",X"05",X"89",X"86",X"10",X"08",X"86",X"8A",X"3C",X"75",X"10",X"03",X"85",
		X"7E",X"90",X"7B",X"7C",X"76",X"91",X"83",X"92",X"9A",X"92",X"96",X"84",X"9E",X"92",X"96",X"96",
		X"92",X"9A",X"92",X"96",X"96",X"9E",X"38",X"3C",X"75",X"10",X"03",X"9C",X"8E",X"7A",X"78",X"78",
		X"7E",X"93",X"9F",X"99",X"94",X"94",X"97",X"94",X"97",X"94",X"99",X"97",X"94",X"97",X"94",X"94",
		X"94",X"97",X"97",X"3C",X"75",X"10",X"02",X"88",X"7E",X"7A",X"78",X"7A",X"7A",X"8E",X"93",X"64",
		X"95",X"95",X"95",X"95",X"98",X"98",X"95",X"98",X"95",X"95",X"98",X"95",X"98",X"98",X"98",X"95",
		X"3C",X"75",X"10",X"03",X"E6",X"E7",X"57",X"72",X"67",X"72",X"4C",X"55",X"55",X"67",X"72",X"4C",
		X"55",X"67",X"72",X"4C",X"55",X"67",X"72",X"4C",X"4C",X"55",X"5F",X"62",X"3C",X"75",X"10",X"03",
		X"E4",X"E5",X"57",X"72",X"6B",X"73",X"73",X"68",X"68",X"6B",X"73",X"73",X"68",X"6B",X"73",X"73",
		X"68",X"6B",X"73",X"73",X"68",X"68",X"5D",X"5D",X"3C",X"75",X"10",X"03",X"E6",X"E7",X"57",X"67",
		X"6A",X"39",X"39",X"67",X"67",X"6A",X"39",X"39",X"67",X"6A",X"39",X"39",X"67",X"6A",X"39",X"39",
		X"67",X"67",X"41",X"65",X"3C",X"75",X"10",X"03",X"A8",X"A9",X"A2",X"A1",X"69",X"3A",X"3A",X"66",
		X"65",X"69",X"3A",X"3A",X"66",X"69",X"3A",X"3A",X"66",X"69",X"3A",X"3A",X"66",X"65",X"69",X"69",
		X"3C",X"75",X"10",X"03",X"AA",X"AB",X"10",X"16",X"3C",X"75",X"10",X"03",X"AF",X"37",X"37",X"37",
		X"37",X"37",X"37",X"37",X"37",X"37",X"37",X"37",X"37",X"37",X"37",X"37",X"37",X"35",X"10",X"06",
		X"3C",X"75",X"10",X"03",X"C4",X"C2",X"10",X"16",X"3C",X"75",X"10",X"03",X"57",X"61",X"10",X"16",
		X"3C",X"75",X"10",X"03",X"57",X"60",X"10",X"16",X"3C",X"75",X"10",X"03",X"57",X"60",X"10",X"16",
		X"3C",X"75",X"10",X"03",X"57",X"41",X"C2",X"10",X"14",X"2F",X"3C",X"75",X"10",X"03",X"57",X"5E",
		X"61",X"10",X"14",X"2F",X"3C",X"75",X"10",X"03",X"57",X"5E",X"62",X"10",X"15",X"3C",X"75",X"10",
		X"03",X"57",X"5D",X"62",X"10",X"15",X"3C",X"75",X"10",X"03",X"57",X"5F",X"62",X"10",X"14",X"2F",
		X"3C",X"75",X"10",X"03",X"57",X"5D",X"61",X"10",X"14",X"2F",X"3C",X"75",X"10",X"03",X"57",X"5E",
		X"60",X"10",X"15",X"3C",X"75",X"10",X"03",X"57",X"5F",X"60",X"10",X"15",X"3C",X"75",X"10",X"03",
		X"57",X"5F",X"61",X"10",X"14",X"2F",X"3C",X"75",X"10",X"03",X"57",X"5E",X"61",X"10",X"14",X"2F",
		X"3C",X"75",X"10",X"03",X"57",X"5D",X"60",X"10",X"15",X"3C",X"75",X"10",X"03",X"57",X"41",X"41",
		X"5A",X"10",X"14",X"3C",X"75",X"10",X"03",X"57",X"5B",X"41",X"61",X"10",X"14",X"3C",X"75",X"10",
		X"03",X"57",X"5B",X"5B",X"41",X"10",X"14",X"3C",X"75",X"10",X"03",X"57",X"41",X"4B",X"4A",X"59",
		X"10",X"10",X"A3",X"A3",X"A3",X"3C",X"75",X"10",X"03",X"57",X"41",X"4B",X"4A",X"41",X"50",X"52",
		X"10",X"02",X"50",X"50",X"50",X"4E",X"4E",X"50",X"50",X"50",X"10",X"02",X"52",X"50",X"6C",X"D0",
		X"D1",X"3C",X"75",X"10",X"03",X"57",X"41",X"56",X"56",X"41",X"59",X"56",X"49",X"48",X"4A",X"4B",
		X"4C",X"4D",X"4D",X"4C",X"4B",X"4A",X"49",X"48",X"56",X"59",X"6E",X"D2",X"D3",X"3C",X"75",X"10",
		X"03",X"57",X"67",X"67",X"41",X"56",X"67",X"67",X"41",X"49",X"44",X"44",X"45",X"56",X"56",X"45",
		X"44",X"44",X"49",X"41",X"67",X"67",X"70",X"D0",X"D1",X"3C",X"75",X"3A",X"07",X"89",X"CB",X"47",
		X"C8",X"3A",X"02",X"89",X"32",X"43",X"8D",X"32",X"34",X"89",X"A7",X"20",X"0F",X"21",X"E3",X"86",
		X"22",X"32",X"89",X"2E",X"82",X"11",X"54",X"27",X"CD",X"07",X"33",X"C9",X"47",X"21",X"A3",X"86",
		X"22",X"32",X"89",X"2E",X"C3",X"11",X"DF",X"FF",X"36",X"DA",X"23",X"36",X"DB",X"19",X"36",X"D8",
		X"23",X"36",X"D9",X"19",X"10",X"F2",X"1E",X"BF",X"19",X"11",X"54",X"27",X"CD",X"07",X"33",X"C9",
		X"10",X"1D",X"10",X"08",X"40",X"10",X"04",X"40",X"10",X"03",X"40",X"10",X"03",X"40",X"00",X"80",
		X"10",X"05",X"10",X"1D",X"10",X"17",X"80",X"80",X"10",X"04",X"10",X"18",X"80",X"10",X"04",X"10",
		X"1D",X"10",X"03",X"40",X"10",X"19",X"10",X"03",X"40",X"10",X"19",X"10",X"1D",X"10",X"04",X"80",
		X"80",X"10",X"17",X"10",X"1A",X"07",X"10",X"02",X"10",X"05",X"80",X"10",X"17",X"10",X"1D",X"10",
		X"1D",X"10",X"05",X"80",X"10",X"14",X"0E",X"10",X"02",X"10",X"1D",X"10",X"03",X"80",X"10",X"19",
		X"FF",X"C2",X"82",X"02",X"10",X"04",X"40",X"10",X"18",X"10",X"1D",X"10",X"1D",X"10",X"04",X"80",
		X"10",X"18",X"10",X"04",X"80",X"10",X"02",X"80",X"10",X"11",X"40",X"10",X"03",X"10",X"07",X"80",
		X"10",X"0B",X"40",X"10",X"05",X"40",X"00",X"10",X"02",X"10",X"08",X"40",X"10",X"04",X"40",X"02",
		X"40",X"10",X"06",X"40",X"10",X"06",X"10",X"02",X"C0",X"10",X"04",X"80",X"40",X"80",X"00",X"00",
		X"00",X"40",X"10",X"02",X"40",X"10",X"02",X"40",X"10",X"02",X"40",X"10",X"03",X"40",X"10",X"02",
		X"FF",X"A2",X"80",X"02",X"10",X"10",X"80",X"80",X"10",X"0B",X"10",X"11",X"80",X"10",X"0B",X"10",
		X"1D",X"10",X"13",X"07",X"10",X"09",X"10",X"13",X"07",X"10",X"09",X"FF",X"A2",X"82",X"0A",X"10",
		X"13",X"0E",X"10",X"09",X"10",X"1D",X"10",X"1D",X"10",X"13",X"0E",X"10",X"09",X"10",X"1D",X"10",
		X"1D",X"10",X"13",X"07",X"10",X"09",X"10",X"13",X"07",X"10",X"09",X"10",X"13",X"0E",X"10",X"09",
		X"FF",X"A2",X"80",X"02",X"10",X"10",X"80",X"80",X"10",X"0B",X"10",X"11",X"80",X"10",X"0B",X"FF",
		X"42",X"81",X"02",X"10",X"13",X"07",X"10",X"09",X"FF",X"C2",X"81",X"02",X"10",X"13",X"0E",X"10",
		X"09",X"FF",X"C2",X"83",X"0E",X"10",X"1D",X"10",X"06",X"07",X"10",X"05",X"40",X"10",X"10",X"10",
		X"1D",X"10",X"10",X"80",X"80",X"10",X"0B",X"10",X"11",X"80",X"10",X"0B",X"10",X"1D",X"10",X"1D",
		X"10",X"13",X"0E",X"10",X"09",X"10",X"01",X"C0",X"C0",X"10",X"1A",X"10",X"01",X"00",X"00",X"10",
		X"1A",X"10",X"01",X"85",X"82",X"10",X"10",X"0E",X"10",X"09",X"10",X"01",X"05",X"02",X"10",X"1A",
		X"10",X"01",X"80",X"80",X"10",X"1A",X"10",X"01",X"00",X"00",X"10",X"04",X"40",X"10",X"15",X"10",
		X"01",X"8D",X"CD",X"10",X"04",X"40",X"10",X"15",X"10",X"01",X"0D",X"4D",X"10",X"1A",X"10",X"01",
		X"83",X"C3",X"10",X"05",X"80",X"80",X"10",X"13",X"10",X"01",X"03",X"43",X"10",X"1A",X"10",X"01",
		X"80",X"C0",X"10",X"06",X"80",X"10",X"13",X"10",X"01",X"00",X"00",X"10",X"05",X"80",X"10",X"14",
		X"FF",X"42",X"83",X"03",X"10",X"08",X"80",X"10",X"09",X"40",X"10",X"0A",X"10",X"0A",X"80",X"10",
		X"07",X"40",X"00",X"10",X"09",X"10",X"1D",X"10",X"09",X"80",X"40",X"00",X"82",X"00",X"40",X"00",
		X"40",X"00",X"00",X"40",X"10",X"09",X"10",X"1D",X"10",X"08",X"40",X"10",X"04",X"40",X"10",X"03",
		X"40",X"10",X"03",X"04",X"10",X"07",X"10",X"1D",X"10",X"05",X"10",X"18",X"10",X"1D",X"10",X"1D",
		X"10",X"03",X"80",X"40",X"10",X"18",X"FF",X"82",X"81",X"02",X"10",X"05",X"40",X"10",X"14",X"8A",
		X"10",X"02",X"10",X"04",X"10",X"16",X"0A",X"10",X"02",X"10",X"1D",X"10",X"05",X"10",X"18",X"10",
		X"04",X"40",X"10",X"15",X"85",X"10",X"02",X"10",X"1A",X"05",X"10",X"02",X"10",X"04",X"80",X"10",
		X"18",X"10",X"04",X"80",X"80",X"10",X"17",X"10",X"05",X"80",X"10",X"14",X"86",X"10",X"02",X"10",
		X"1A",X"06",X"10",X"02",X"10",X"1D",X"10",X"1D",X"10",X"04",X"80",X"80",X"10",X"17",X"10",X"06",
		X"80",X"10",X"16",X"10",X"05",X"80",X"80",X"10",X"16",X"10",X"08",X"40",X"40",X"10",X"02",X"40",
		X"40",X"40",X"40",X"10",X"0D",X"10",X"06",X"40",X"00",X"40",X"40",X"10",X"02",X"40",X"40",X"40",
		X"40",X"10",X"0D",X"10",X"04",X"40",X"10",X"03",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",
		X"10",X"0D",X"10",X"03",X"E6",X"E7",X"8E",X"7A",X"7E",X"93",X"64",X"95",X"95",X"98",X"95",X"95",
		X"98",X"98",X"95",X"98",X"95",X"95",X"98",X"95",X"98",X"98",X"98",X"95",X"3C",X"75",X"10",X"03",
		X"E4",X"E5",X"7E",X"7B",X"79",X"93",X"9F",X"99",X"99",X"94",X"94",X"97",X"94",X"97",X"94",X"99",
		X"97",X"94",X"97",X"94",X"94",X"94",X"97",X"97",X"3C",X"75",X"10",X"03",X"E6",X"E7",X"9C",X"79",
		X"79",X"91",X"83",X"92",X"92",X"9A",X"92",X"96",X"84",X"9E",X"92",X"96",X"96",X"92",X"9A",X"92",
		X"96",X"96",X"9E",X"38",X"3C",X"75",X"10",X"03",X"A8",X"A9",X"9B",X"7E",X"88",X"10",X"07",X"89",
		X"86",X"10",X"08",X"86",X"8A",X"3C",X"75",X"10",X"03",X"AA",X"AB",X"87",X"8C",X"10",X"13",X"8B",
		X"3C",X"75",X"10",X"03",X"AF",X"37",X"37",X"37",X"34",X"10",X"13",X"3C",X"75",X"10",X"1B",X"3C",
		X"75",X"10",X"1B",X"3C",X"75",X"10",X"1B",X"3C",X"75",X"10",X"1B",X"3C",X"75",X"10",X"1B",X"3C",
		X"75",X"10",X"1B",X"3C",X"75",X"10",X"1B",X"3C",X"75",X"10",X"1B",X"3C",X"75",X"10",X"1B",X"3C",
		X"75",X"10",X"1B",X"3C",X"75",X"10",X"1B",X"3C",X"75",X"10",X"1B",X"3C",X"75",X"10",X"1B",X"3C",
		X"75",X"87",X"87",X"10",X"19",X"3C",X"75",X"9C",X"7E",X"87",X"10",X"18",X"3C",X"75",X"85",X"76",
		X"76",X"87",X"10",X"17",X"3C",X"75",X"7E",X"7B",X"90",X"8F",X"8C",X"10",X"16",X"3C",X"75",X"7F",
		X"7B",X"7C",X"76",X"76",X"87",X"10",X"14",X"8B",X"3C",X"75",X"85",X"79",X"76",X"76",X"79",X"76",
		X"88",X"10",X"12",X"86",X"8A",X"3C",X"75",X"85",X"7E",X"90",X"7B",X"7C",X"76",X"91",X"83",X"39",
		X"39",X"39",X"39",X"39",X"39",X"39",X"39",X"39",X"39",X"39",X"39",X"39",X"39",X"39",X"39",X"39",
		X"9E",X"38",X"3C",X"75",X"85",X"8E",X"7A",X"78",X"78",X"7E",X"93",X"9F",X"3A",X"3A",X"3A",X"3A",
		X"3A",X"3A",X"3A",X"3A",X"3A",X"3A",X"3A",X"3A",X"3A",X"3A",X"3A",X"3A",X"3A",X"97",X"94",X"3C",
		X"75",X"7E",X"7A",X"78",X"7A",X"7A",X"8E",X"93",X"64",X"95",X"98",X"95",X"95",X"98",X"98",X"95",
		X"98",X"98",X"95",X"98",X"95",X"95",X"98",X"95",X"98",X"98",X"98",X"95",X"3C",X"75",X"10",X"05",
		X"80",X"80",X"C0",X"00",X"00",X"80",X"80",X"C0",X"C0",X"80",X"80",X"C0",X"80",X"80",X"C0",X"80",
		X"80",X"C0",X"80",X"80",X"80",X"C0",X"00",X"00",X"10",X"05",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"C0",X"82",X"C0",X"80",X"80",X"80",X"80",X"80",X"80",X"C0",X"80",X"80",X"80",X"80",
		X"00",X"00",X"10",X"05",X"00",X"00",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"C0",X"80",X"80",X"80",X"80",X"80",X"C0",X"00",X"10",X"02",X"10",X"05",X"40",X"00",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"C0",X"80",X"00",X"00",X"10",X"05",X"C0",X"80",X"10",X"13",X"80",X"00",X"00",X"FF",
		X"A2",X"82",X"0D",X"40",X"10",X"1C",X"10",X"01",X"80",X"10",X"1B",X"10",X"1D",X"10",X"1D",X"00",
		X"80",X"10",X"1B",X"00",X"80",X"10",X"02",X"80",X"10",X"14",X"40",X"10",X"03",X"10",X"04",X"80",
		X"10",X"14",X"40",X"10",X"03",X"10",X"05",X"40",X"10",X"17",X"10",X"04",X"80",X"40",X"80",X"00",
		X"00",X"40",X"40",X"10",X"02",X"40",X"10",X"02",X"40",X"10",X"02",X"40",X"10",X"03",X"40",X"10",
		X"05",X"10",X"03",X"E6",X"E7",X"57",X"72",X"67",X"72",X"4C",X"55",X"55",X"67",X"72",X"4C",X"55",
		X"67",X"72",X"4C",X"55",X"67",X"72",X"4C",X"63",X"31",X"4F",X"4F",X"3C",X"75",X"10",X"03",X"E4",
		X"E5",X"57",X"72",X"6B",X"73",X"73",X"68",X"68",X"6B",X"73",X"73",X"68",X"6B",X"73",X"73",X"68",
		X"6B",X"73",X"73",X"2E",X"30",X"3D",X"81",X"3C",X"75",X"10",X"03",X"E6",X"E7",X"57",X"67",X"6A",
		X"39",X"39",X"67",X"67",X"6A",X"39",X"39",X"67",X"6A",X"39",X"39",X"67",X"6A",X"39",X"39",X"2E",
		X"32",X"42",X"BD",X"3C",X"75",X"10",X"03",X"A8",X"A9",X"A2",X"A1",X"69",X"3A",X"3A",X"66",X"65",
		X"69",X"3A",X"3A",X"66",X"69",X"3A",X"3A",X"66",X"69",X"3A",X"3A",X"2E",X"32",X"3D",X"81",X"3C",
		X"75",X"10",X"03",X"AA",X"AB",X"10",X"12",X"33",X"30",X"42",X"BD",X"3C",X"75",X"10",X"03",X"AF",
		X"37",X"37",X"37",X"34",X"10",X"10",X"6D",X"58",X"58",X"3C",X"75",X"10",X"03",X"87",X"87",X"10",
		X"16",X"3C",X"75",X"10",X"03",X"9B",X"9D",X"88",X"10",X"15",X"3C",X"75",X"10",X"03",X"9C",X"82",
		X"88",X"10",X"15",X"3C",X"75",X"10",X"03",X"79",X"79",X"88",X"10",X"01",X"00",X"10",X"13",X"3C",
		X"75",X"10",X"03",X"9C",X"82",X"87",X"10",X"01",X"00",X"10",X"12",X"2F",X"3C",X"75",X"10",X"03",
		X"85",X"76",X"87",X"10",X"14",X"2F",X"3C",X"75",X"10",X"03",X"9C",X"76",X"87",X"10",X"15",X"3C",
		X"75",X"10",X"03",X"9C",X"79",X"9B",X"10",X"15",X"3C",X"75",X"10",X"03",X"79",X"76",X"87",X"10",
		X"14",X"2F",X"3C",X"75",X"10",X"03",X"80",X"8D",X"10",X"02",X"24",X"10",X"12",X"2F",X"3C",X"75",
		X"10",X"03",X"80",X"76",X"87",X"10",X"01",X"1E",X"10",X"13",X"3C",X"75",X"10",X"03",X"85",X"76",
		X"9B",X"10",X"01",X"19",X"10",X"13",X"3C",X"75",X"10",X"03",X"85",X"82",X"9B",X"10",X"01",X"1F",
		X"10",X"12",X"2F",X"3C",X"75",X"10",X"03",X"9C",X"79",X"9B",X"10",X"01",X"20",X"10",X"12",X"2F",
		X"3C",X"75",X"10",X"03",X"9C",X"79",X"9D",X"88",X"10",X"14",X"3C",X"75",X"10",X"03",X"85",X"76",
		X"76",X"87",X"10",X"14",X"3C",X"75",X"10",X"03",X"7E",X"7B",X"90",X"8F",X"8C",X"10",X"13",X"3C",
		X"75",X"B7",X"B8",X"B9",X"7F",X"7B",X"7C",X"76",X"76",X"87",X"10",X"11",X"8B",X"3C",X"75",X"B6",
		X"B1",X"B6",X"85",X"79",X"76",X"76",X"79",X"9D",X"88",X"10",X"05",X"89",X"86",X"10",X"08",X"86",
		X"8A",X"3C",X"75",X"B4",X"B5",X"B4",X"85",X"7E",X"90",X"7B",X"7C",X"76",X"91",X"83",X"92",X"9A",
		X"92",X"96",X"84",X"9E",X"92",X"96",X"96",X"92",X"9A",X"92",X"96",X"96",X"9E",X"38",X"3C",X"75",
		X"10",X"03",X"9C",X"8E",X"7A",X"78",X"78",X"7E",X"93",X"9F",X"99",X"94",X"94",X"97",X"94",X"97",
		X"94",X"99",X"97",X"94",X"97",X"94",X"94",X"94",X"97",X"97",X"3C",X"75",X"10",X"02",X"88",X"7E",
		X"7A",X"78",X"7A",X"7A",X"8E",X"93",X"64",X"95",X"95",X"95",X"95",X"98",X"98",X"95",X"98",X"95",
		X"95",X"98",X"95",X"98",X"98",X"98",X"95",X"3C",X"75",X"10",X"1D",X"10",X"08",X"40",X"10",X"04",
		X"40",X"10",X"03",X"40",X"10",X"03",X"40",X"00",X"80",X"10",X"05",X"10",X"1D",X"10",X"17",X"80",
		X"80",X"10",X"04",X"10",X"18",X"80",X"10",X"04",X"10",X"1D",X"10",X"03",X"40",X"10",X"19",X"10",
		X"03",X"40",X"10",X"19",X"10",X"1D",X"10",X"04",X"80",X"80",X"10",X"17",X"10",X"1A",X"8A",X"10",
		X"02",X"10",X"05",X"80",X"10",X"14",X"0A",X"10",X"02",X"10",X"1D",X"10",X"1D",X"10",X"05",X"80",
		X"10",X"14",X"85",X"10",X"02",X"10",X"1A",X"05",X"10",X"02",X"10",X"03",X"80",X"10",X"19",X"10",
		X"1D",X"10",X"1A",X"86",X"10",X"02",X"10",X"1A",X"06",X"10",X"02",X"10",X"04",X"40",X"10",X"18",
		X"10",X"1D",X"10",X"1D",X"80",X"80",X"80",X"00",X"80",X"10",X"18",X"80",X"00",X"C0",X"00",X"80",
		X"10",X"02",X"80",X"10",X"11",X"40",X"10",X"03",X"80",X"80",X"C0",X"10",X"04",X"80",X"10",X"0B",
		X"40",X"10",X"05",X"40",X"00",X"10",X"02",X"10",X"02",X"C0",X"10",X"05",X"40",X"10",X"04",X"40",
		X"02",X"40",X"10",X"06",X"40",X"10",X"06",X"10",X"02",X"C0",X"10",X"04",X"80",X"40",X"80",X"00",
		X"00",X"00",X"40",X"10",X"02",X"40",X"10",X"02",X"40",X"10",X"02",X"40",X"10",X"03",X"40",X"10",
		X"02",X"3A",X"FB",X"89",X"A7",X"20",X"22",X"21",X"C5",X"6A",X"11",X"00",X"00",X"7E",X"FE",X"C9",
		X"28",X"08",X"83",X"5F",X"30",X"01",X"14",X"23",X"18",X"F3",X"21",X"19",X"51",X"7B",X"BE",X"C3",
		X"C5",X"6A",X"7A",X"23",X"BE",X"C2",X"2C",X"46",X"C9",X"ED",X"1B",X"3A",X"07",X"89",X"CB",X"47",
		X"28",X"1F",X"CD",X"C5",X"54",X"CD",X"19",X"55",X"CD",X"64",X"55",X"3A",X"61",X"8F",X"A7",X"28",
		X"04",X"CD",X"71",X"11",X"C9",X"CD",X"46",X"51",X"3A",X"6D",X"8D",X"A7",X"C0",X"CD",X"E8",X"56",
		X"C9",X"CD",X"B0",X"53",X"18",X"EF",X"CD",X"50",X"51",X"CD",X"F6",X"52",X"CD",X"34",X"53",X"C9",
		X"3A",X"6D",X"8D",X"A7",X"C0",X"21",X"9A",X"51",X"3A",X"07",X"89",X"E6",X"0F",X"CD",X"45",X"0C",
		X"EB",X"3A",X"01",X"89",X"FE",X"07",X"D8",X"BE",X"28",X"05",X"D0",X"23",X"23",X"18",X"F8",X"32",
		X"6D",X"8D",X"23",X"7E",X"47",X"32",X"74",X"8D",X"21",X"64",X"52",X"CD",X"45",X"0C",X"1A",X"32",
		X"73",X"8D",X"13",X"ED",X"53",X"71",X"8D",X"78",X"21",X"B0",X"52",X"CD",X"45",X"0C",X"ED",X"53",
		X"6F",X"8D",X"AF",X"32",X"7B",X"8D",X"32",X"7E",X"8D",X"C9",X"BA",X"51",X"C2",X"51",X"CA",X"51",
		X"D4",X"51",X"DE",X"51",X"E8",X"51",X"F4",X"51",X"00",X"52",X"0C",X"52",X"16",X"52",X"20",X"52",
		X"2A",X"52",X"36",X"52",X"42",X"52",X"4E",X"52",X"5A",X"52",X"20",X"00",X"18",X"00",X"10",X"00",
		X"05",X"02",X"20",X"04",X"18",X"02",X"10",X"05",X"05",X"02",X"28",X"05",X"20",X"00",X"18",X"05",
		X"10",X"01",X"05",X"04",X"28",X"01",X"20",X"02",X"18",X"02",X"10",X"01",X"05",X"04",X"28",X"02",
		X"20",X"01",X"18",X"03",X"10",X"04",X"05",X"04",X"30",X"00",X"28",X"06",X"20",X"05",X"18",X"03",
		X"10",X"00",X"05",X"04",X"30",X"08",X"28",X"04",X"20",X"05",X"18",X"06",X"10",X"07",X"05",X"04",
		X"30",X"06",X"28",X"07",X"20",X"00",X"18",X"05",X"10",X"02",X"05",X"04",X"28",X"09",X"20",X"00",
		X"18",X"05",X"10",X"03",X"05",X"04",X"28",X"01",X"20",X"02",X"18",X"02",X"10",X"07",X"05",X"04",
		X"28",X"02",X"20",X"01",X"18",X"03",X"10",X"08",X"05",X"04",X"30",X"04",X"28",X"07",X"20",X"02",
		X"18",X"06",X"10",X"01",X"05",X"04",X"30",X"04",X"28",X"01",X"20",X"06",X"18",X"00",X"10",X"09",
		X"05",X"04",X"30",X"07",X"28",X"06",X"20",X"00",X"18",X"05",X"10",X"02",X"05",X"04",X"2B",X"09",
		X"24",X"08",X"1C",X"04",X"14",X"07",X"0D",X"02",X"05",X"02",X"28",X"00",X"20",X"02",X"18",X"06",
		X"10",X"07",X"05",X"04",X"78",X"52",X"7F",X"52",X"86",X"52",X"8D",X"52",X"94",X"52",X"9B",X"52",
		X"9B",X"52",X"9B",X"52",X"A2",X"52",X"A9",X"52",X"01",X"1E",X"18",X"14",X"10",X"10",X"FF",X"01",
		X"30",X"30",X"34",X"30",X"30",X"FF",X"01",X"18",X"50",X"38",X"38",X"30",X"FF",X"01",X"38",X"38",
		X"58",X"18",X"30",X"FF",X"01",X"38",X"38",X"38",X"38",X"38",X"FF",X"01",X"30",X"30",X"30",X"30",
		X"30",X"FF",X"01",X"50",X"20",X"3E",X"60",X"40",X"FF",X"01",X"10",X"60",X"58",X"60",X"30",X"FF",
		X"C4",X"52",X"C9",X"52",X"CE",X"52",X"D3",X"52",X"D8",X"52",X"DD",X"52",X"E2",X"52",X"E7",X"52",
		X"EC",X"52",X"F1",X"52",X"08",X"0A",X"0D",X"10",X"12",X"13",X"10",X"0D",X"0A",X"07",X"0E",X"10",
		X"0B",X"09",X"07",X"10",X"0E",X"0C",X"08",X"0A",X"10",X"0E",X"0C",X"0A",X"08",X"08",X"08",X"08",
		X"08",X"08",X"0D",X"0D",X"0D",X"0D",X"0D",X"10",X"10",X"10",X"10",X"10",X"14",X"08",X"0E",X"14",
		X"08",X"0E",X"14",X"07",X"14",X"07",X"3A",X"6D",X"8D",X"A7",X"C8",X"3A",X"6E",X"8D",X"A7",X"C0",
		X"01",X"00",X"06",X"21",X"E0",X"8A",X"11",X"17",X"00",X"7E",X"2C",X"B6",X"20",X"01",X"0C",X"19",
		X"10",X"F7",X"79",X"FE",X"04",X"D8",X"32",X"6E",X"8D",X"11",X"F3",X"0B",X"06",X"17",X"AF",X"6F",
		X"67",X"1A",X"E7",X"1B",X"10",X"FB",X"3E",X"EB",X"85",X"20",X"04",X"7C",X"C6",X"F7",X"C8",X"21",
		X"E8",X"89",X"34",X"C9",X"3A",X"6E",X"8D",X"A7",X"C8",X"ED",X"5B",X"71",X"8D",X"1A",X"3C",X"20",
		X"14",X"3A",X"6D",X"8D",X"47",X"3A",X"01",X"89",X"B8",X"D0",X"AF",X"32",X"6D",X"8D",X"32",X"6E",
		X"8D",X"32",X"07",X"8D",X"C9",X"21",X"73",X"8D",X"35",X"C0",X"3D",X"77",X"13",X"ED",X"53",X"71",
		X"8D",X"DD",X"21",X"E0",X"8A",X"11",X"18",X"00",X"06",X"06",X"D9",X"CD",X"74",X"53",X"D9",X"DD",
		X"19",X"10",X"F7",X"C9",X"DD",X"7E",X"00",X"DD",X"B6",X"01",X"C0",X"21",X"79",X"8D",X"34",X"DD",
		X"36",X"00",X"01",X"3A",X"07",X"89",X"1E",X"1D",X"CB",X"47",X"20",X"02",X"1E",X"04",X"CD",X"A0",
		X"53",X"21",X"A6",X"53",X"3A",X"74",X"8D",X"E7",X"DD",X"B6",X"07",X"DD",X"77",X"07",X"F1",X"C9",
		X"0E",X"FF",X"CD",X"33",X"57",X"C9",X"14",X"24",X"34",X"44",X"54",X"64",X"74",X"84",X"94",X"A4",
		X"A7",X"C8",X"3A",X"59",X"8D",X"A7",X"C0",X"3A",X"5F",X"8A",X"A7",X"C0",X"3C",X"32",X"59",X"8D",
		X"DD",X"21",X"30",X"8C",X"21",X"02",X"59",X"E7",X"DD",X"77",X"09",X"ED",X"44",X"DD",X"77",X"0A",
		X"DD",X"36",X"00",X"01",X"DD",X"36",X"02",X"0B",X"AF",X"DD",X"77",X"03",X"DD",X"36",X"04",X"04",
		X"DD",X"77",X"05",X"DD",X"77",X"06",X"2F",X"32",X"4B",X"8D",X"11",X"03",X"42",X"CD",X"1E",X"38",
		X"3A",X"07",X"89",X"CB",X"3F",X"3C",X"FE",X"07",X"38",X"02",X"3E",X"06",X"32",X"5C",X"8D",X"21",
		X"07",X"54",X"E7",X"32",X"5D",X"8D",X"C9",X"FF",X"20",X"18",X"0C",X"0C",X"0B",X"3A",X"07",X"89",
		X"E6",X"01",X"C8",X"AF",X"21",X"01",X"8D",X"06",X"06",X"D7",X"21",X"11",X"8D",X"06",X"06",X"D7",
		X"DD",X"21",X"30",X"8C",X"11",X"18",X"00",X"06",X"03",X"D9",X"CD",X"33",X"54",X"D9",X"DD",X"19",
		X"10",X"F7",X"C9",X"DD",X"7E",X"00",X"DD",X"B6",X"01",X"C0",X"DD",X"36",X"00",X"01",X"AF",X"DD",
		X"77",X"02",X"DD",X"77",X"05",X"DD",X"36",X"03",X"60",X"DD",X"36",X"04",X"1B",X"DD",X"77",X"0E",
		X"21",X"D4",X"55",X"3A",X"01",X"8D",X"4F",X"E7",X"DD",X"77",X"06",X"21",X"D7",X"55",X"79",X"E7",
		X"ED",X"44",X"DD",X"77",X"0A",X"21",X"1F",X"56",X"79",X"CD",X"45",X"0C",X"1A",X"DD",X"77",X"17",
		X"21",X"57",X"56",X"CD",X"45",X"0C",X"DD",X"73",X"0C",X"DD",X"72",X"0D",X"DD",X"36",X"11",X"40",
		X"CD",X"06",X"40",X"79",X"3C",X"32",X"01",X"8D",X"C9",X"DD",X"36",X"00",X"01",X"AF",X"DD",X"77",
		X"02",X"DD",X"77",X"05",X"DD",X"36",X"03",X"60",X"DD",X"36",X"04",X"1B",X"DD",X"70",X"06",X"DD",
		X"7E",X"17",X"4F",X"21",X"57",X"56",X"CD",X"45",X"0C",X"CD",X"1E",X"38",X"DD",X"36",X"11",X"40",
		X"79",X"21",X"D7",X"55",X"E7",X"3A",X"07",X"89",X"E6",X"07",X"4F",X"87",X"81",X"E7",X"ED",X"44",
		X"DD",X"77",X"0A",X"F1",X"C9",X"3A",X"07",X"89",X"FE",X"04",X"30",X"0F",X"FE",X"02",X"3A",X"20",
		X"88",X"38",X"05",X"FE",X"02",X"D8",X"18",X"03",X"FE",X"03",X"D8",X"21",X"04",X"8D",X"35",X"C0",
		X"21",X"EF",X"55",X"3A",X"12",X"8D",X"E6",X"0F",X"E7",X"32",X"04",X"8D",X"21",X"12",X"8D",X"34",
		X"DD",X"21",X"30",X"8C",X"11",X"18",X"00",X"06",X"01",X"D9",X"DD",X"7E",X"00",X"DD",X"B6",X"01",
		X"20",X"11",X"06",X"0B",X"21",X"37",X"56",X"3A",X"12",X"8D",X"E6",X"0F",X"E7",X"DD",X"77",X"17",
		X"CD",X"89",X"54",X"D9",X"DD",X"19",X"10",X"E1",X"C9",X"3A",X"07",X"89",X"FE",X"02",X"30",X"06",
		X"3A",X"20",X"88",X"FE",X"02",X"D8",X"21",X"05",X"8D",X"35",X"C0",X"21",X"FF",X"55",X"3A",X"13",
		X"8D",X"E6",X"0F",X"E7",X"32",X"05",X"8D",X"21",X"13",X"8D",X"34",X"DD",X"21",X"48",X"8C",X"11",
		X"18",X"00",X"06",X"01",X"D9",X"DD",X"7E",X"00",X"DD",X"B6",X"01",X"20",X"11",X"06",X"0F",X"21",
		X"47",X"56",X"3A",X"13",X"8D",X"E6",X"0F",X"E7",X"DD",X"77",X"17",X"CD",X"89",X"54",X"D9",X"DD",
		X"19",X"10",X"E1",X"C9",X"21",X"06",X"8D",X"35",X"C0",X"21",X"0F",X"56",X"3A",X"14",X"8D",X"E6",
		X"0F",X"E7",X"32",X"06",X"8D",X"21",X"14",X"8D",X"34",X"DD",X"21",X"60",X"8C",X"11",X"18",X"00",
		X"3A",X"07",X"89",X"FE",X"04",X"30",X"0B",X"3A",X"20",X"88",X"A7",X"C8",X"FE",X"04",X"06",X"01",
		X"38",X"02",X"06",X"02",X"D9",X"DD",X"7E",X"00",X"DD",X"B6",X"01",X"20",X"31",X"11",X"AD",X"0B",
		X"21",X"B5",X"55",X"06",X"08",X"1A",X"86",X"20",X"06",X"13",X"23",X"10",X"F8",X"18",X"0E",X"21",
		X"1E",X"88",X"34",X"18",X"08",X"AA",X"7A",X"AD",X"7A",X"B2",X"7A",X"B5",X"7A",X"06",X"13",X"21",
		X"27",X"56",X"3A",X"14",X"8D",X"E6",X"0F",X"E7",X"DD",X"77",X"17",X"CD",X"89",X"54",X"D9",X"DD",
		X"19",X"10",X"C1",X"C9",X"0B",X"0F",X"13",X"10",X"18",X"20",X"20",X"18",X"10",X"28",X"18",X"20",
		X"10",X"18",X"20",X"18",X"20",X"10",X"28",X"18",X"20",X"10",X"18",X"28",X"18",X"18",X"20",X"40",
		X"50",X"60",X"70",X"80",X"90",X"A0",X"B0",X"C0",X"D0",X"E0",X"F0",X"10",X"20",X"30",X"40",X"F0",
		X"E0",X"D0",X"C0",X"B0",X"A0",X"90",X"80",X"70",X"60",X"50",X"40",X"30",X"20",X"10",X"F0",X"20",
		X"30",X"40",X"20",X"20",X"50",X"40",X"30",X"20",X"60",X"20",X"30",X"40",X"70",X"30",X"40",X"27",
		X"56",X"37",X"56",X"47",X"56",X"47",X"56",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"02",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"03",X"01",X"01",X"01",X"01",X"01",X"00",X"03",
		X"03",X"01",X"01",X"00",X"00",X"01",X"01",X"02",X"02",X"02",X"02",X"02",X"02",X"01",X"02",X"02",
		X"00",X"02",X"03",X"02",X"03",X"03",X"02",X"61",X"56",X"7C",X"56",X"97",X"56",X"B2",X"56",X"CD",
		X"56",X"44",X"3C",X"10",X"44",X"3D",X"10",X"44",X"3E",X"10",X"44",X"E1",X"10",X"44",X"E2",X"10",
		X"44",X"E1",X"10",X"44",X"E2",X"10",X"44",X"E1",X"10",X"FF",X"6D",X"56",X"41",X"3C",X"10",X"41",
		X"3D",X"10",X"41",X"3E",X"10",X"41",X"E1",X"10",X"41",X"E2",X"10",X"41",X"E1",X"10",X"41",X"E2",
		X"10",X"41",X"E1",X"10",X"FF",X"88",X"56",X"49",X"3C",X"10",X"49",X"3D",X"10",X"49",X"3E",X"10",
		X"49",X"E1",X"10",X"49",X"E2",X"10",X"49",X"E1",X"10",X"49",X"E2",X"10",X"49",X"E1",X"10",X"FF",
		X"A3",X"56",X"4C",X"3C",X"10",X"4C",X"3D",X"10",X"4C",X"3E",X"10",X"4C",X"E1",X"10",X"4C",X"E2",
		X"10",X"4C",X"E1",X"10",X"4C",X"E2",X"10",X"4C",X"E1",X"10",X"FF",X"BE",X"56",X"40",X"3C",X"10",
		X"40",X"3D",X"10",X"40",X"3E",X"10",X"40",X"E1",X"10",X"40",X"E2",X"10",X"40",X"E1",X"10",X"40",
		X"E2",X"10",X"40",X"E1",X"10",X"FF",X"D9",X"56",X"3A",X"07",X"8D",X"A7",X"28",X"05",X"3D",X"32",
		X"07",X"8D",X"C9",X"3A",X"07",X"89",X"CB",X"47",X"CA",X"71",X"58",X"3A",X"01",X"89",X"21",X"40",
		X"8D",X"96",X"C8",X"D8",X"4F",X"3A",X"00",X"89",X"FE",X"03",X"38",X"04",X"06",X"06",X"18",X"03",
		X"C6",X"04",X"47",X"3A",X"40",X"8D",X"B8",X"D0",X"DD",X"21",X"E0",X"8A",X"06",X"06",X"1E",X"1D",
		X"CD",X"2B",X"57",X"11",X"18",X"00",X"DD",X"19",X"10",X"F4",X"C9",X"DD",X"7E",X"00",X"DD",X"B6",
		X"01",X"0F",X"D8",X"41",X"DD",X"36",X"00",X"01",X"DD",X"36",X"02",X"03",X"DD",X"73",X"04",X"AF",
		X"DD",X"77",X"03",X"DD",X"77",X"05",X"DD",X"77",X"06",X"DD",X"77",X"08",X"DD",X"36",X"07",X"01",
		X"DD",X"77",X"0B",X"21",X"E0",X"58",X"3A",X"07",X"89",X"E6",X"01",X"20",X"03",X"21",X"02",X"59",
		X"3A",X"20",X"88",X"FE",X"03",X"38",X"02",X"3E",X"03",X"4F",X"3A",X"08",X"89",X"FE",X"04",X"38",
		X"05",X"3A",X"4C",X"8D",X"81",X"4F",X"3A",X"07",X"89",X"CB",X"47",X"CC",X"B4",X"57",X"3A",X"07",
		X"89",X"81",X"4F",X"FE",X"20",X"38",X"02",X"3E",X"1F",X"4F",X"E7",X"DD",X"77",X"09",X"ED",X"44",
		X"DD",X"77",X"0A",X"11",X"29",X"38",X"CD",X"1E",X"38",X"21",X"9B",X"58",X"3A",X"07",X"89",X"E6",
		X"01",X"20",X"03",X"21",X"C0",X"58",X"79",X"E7",X"32",X"07",X"8D",X"21",X"40",X"8D",X"34",X"CD",
		X"C3",X"57",X"F1",X"C9",X"3A",X"01",X"89",X"FE",X"03",X"D0",X"3A",X"7D",X"8D",X"D6",X"0C",X"D8",
		X"81",X"4F",X"C9",X"05",X"28",X"6F",X"21",X"46",X"8D",X"7E",X"A7",X"28",X"2D",X"FE",X"07",X"30",
		X"29",X"34",X"2C",X"7E",X"A7",X"28",X"0A",X"35",X"DD",X"36",X"13",X"02",X"DD",X"36",X"16",X"01",
		X"C9",X"2C",X"7E",X"A7",X"28",X"0A",X"35",X"DD",X"36",X"13",X"01",X"DD",X"36",X"16",X"C1",X"C9",
		X"2C",X"7E",X"A7",X"C8",X"35",X"DD",X"36",X"16",X"41",X"C9",X"36",X"01",X"3A",X"07",X"89",X"CB",
		X"47",X"28",X"25",X"3A",X"00",X"89",X"4F",X"3A",X"4C",X"8D",X"81",X"FE",X"20",X"38",X"02",X"3E",
		X"1F",X"4F",X"EB",X"21",X"22",X"59",X"87",X"81",X"E7",X"13",X"12",X"23",X"13",X"7E",X"12",X"23",
		X"13",X"7E",X"12",X"06",X"FF",X"C3",X"C3",X"57",X"FE",X"20",X"38",X"02",X"3E",X"1F",X"4F",X"EB",
		X"21",X"85",X"59",X"18",X"E1",X"3A",X"4A",X"8D",X"A7",X"20",X"8B",X"3E",X"01",X"32",X"4A",X"8D",
		X"DD",X"77",X"0B",X"DD",X"36",X"13",X"03",X"DD",X"77",X"16",X"DD",X"36",X"07",X"02",X"11",X"47",
		X"38",X"CD",X"1E",X"38",X"21",X"B5",X"0B",X"06",X"52",X"AF",X"57",X"5E",X"83",X"30",X"01",X"14",
		X"23",X"10",X"F8",X"D6",X"C1",X"20",X"04",X"3E",X"1D",X"BA",X"C8",X"3E",X"01",X"32",X"2B",X"88",
		X"C9",X"32",X"00",X"89",X"3A",X"01",X"89",X"21",X"40",X"8D",X"96",X"C8",X"D8",X"3A",X"40",X"8D",
		X"FE",X"06",X"D0",X"3E",X"01",X"32",X"4A",X"8D",X"DD",X"21",X"E0",X"8A",X"06",X"06",X"1E",X"04",
		X"CD",X"2B",X"57",X"11",X"18",X"00",X"DD",X"19",X"10",X"F4",X"C9",X"80",X"80",X"78",X"74",X"70",
		X"6C",X"68",X"60",X"50",X"48",X"40",X"38",X"30",X"2C",X"28",X"24",X"20",X"1E",X"1C",X"1A",X"18",
		X"17",X"17",X"17",X"17",X"16",X"16",X"16",X"16",X"15",X"15",X"15",X"15",X"14",X"14",X"14",X"14",
		X"80",X"70",X"60",X"50",X"48",X"40",X"38",X"30",X"2C",X"28",X"24",X"20",X"1E",X"1C",X"1A",X"18",
		X"17",X"17",X"17",X"17",X"16",X"16",X"16",X"16",X"15",X"15",X"15",X"15",X"14",X"14",X"14",X"14",
		X"10",X"10",X"10",X"10",X"11",X"11",X"12",X"12",X"13",X"13",X"13",X"13",X"14",X"14",X"15",X"15",
		X"15",X"15",X"17",X"17",X"18",X"18",X"19",X"19",X"1A",X"1A",X"1A",X"1A",X"1B",X"1B",X"1B",X"1B",
		X"1C",X"1C",X"10",X"10",X"12",X"12",X"14",X"14",X"15",X"15",X"16",X"16",X"17",X"17",X"18",X"18",
		X"19",X"19",X"19",X"19",X"1A",X"1A",X"1B",X"1B",X"1B",X"1B",X"1C",X"1C",X"1C",X"1C",X"1D",X"1D",
		X"1E",X"1E",X"00",X"00",X"01",X"00",X"00",X"02",X"00",X"00",X"03",X"00",X"00",X"04",X"00",X"00",
		X"05",X"00",X"01",X"03",X"00",X"01",X"04",X"00",X"01",X"05",X"00",X"02",X"02",X"00",X"02",X"03",
		X"00",X"02",X"04",X"00",X"03",X"01",X"00",X"03",X"02",X"00",X"03",X"03",X"00",X"04",X"01",X"00",
		X"04",X"02",X"00",X"05",X"00",X"00",X"05",X"01",X"00",X"06",X"00",X"00",X"05",X"01",X"00",X"06",
		X"00",X"00",X"05",X"01",X"00",X"06",X"00",X"00",X"04",X"02",X"00",X"06",X"00",X"00",X"06",X"00",
		X"00",X"06",X"00",X"00",X"06",X"00",X"00",X"06",X"00",X"00",X"06",X"00",X"00",X"06",X"00",X"00",
		X"06",X"00",X"00",X"06",X"00",X"00",X"00",X"01",X"00",X"00",X"03",X"00",X"00",X"06",X"00",X"01",
		X"04",X"00",X"01",X"05",X"00",X"02",X"03",X"00",X"02",X"04",X"00",X"03",X"01",X"00",X"03",X"02",
		X"00",X"03",X"03",X"00",X"04",X"02",X"00",X"05",X"00",X"00",X"05",X"01",X"01",X"02",X"01",X"01",
		X"01",X"03",X"01",X"01",X"04",X"01",X"02",X"03",X"02",X"00",X"00",X"02",X"01",X"02",X"02",X"00",
		X"01",X"02",X"02",X"01",X"03",X"01",X"01",X"03",X"00",X"01",X"03",X"02",X"00",X"03",X"00",X"02",
		X"03",X"00",X"00",X"03",X"01",X"02",X"03",X"00",X"03",X"04",X"01",X"00",X"04",X"01",X"00",X"04",
		X"00",X"02",X"04",X"00",X"00",X"06",X"00",X"00",X"3A",X"2C",X"88",X"FE",X"0F",X"C8",X"3A",X"2F",
		X"88",X"FE",X"0F",X"C8",X"CD",X"06",X"5A",X"CD",X"56",X"5A",X"CD",X"1F",X"5A",X"CD",X"9C",X"5A",
		X"CD",X"6D",X"7E",X"C3",X"C0",X"5A",X"3A",X"10",X"88",X"0F",X"0F",X"0F",X"21",X"29",X"88",X"CB",
		X"16",X"7E",X"E6",X"07",X"FE",X"01",X"C0",X"CD",X"09",X"0F",X"3E",X"01",X"C3",X"8C",X"5A",X"3A",
		X"10",X"88",X"21",X"2D",X"88",X"0F",X"0F",X"CB",X"16",X"7E",X"E6",X"07",X"FE",X"01",X"C0",X"EB",
		X"CD",X"09",X"0F",X"21",X"26",X"88",X"34",X"EB",X"23",X"7E",X"C6",X"10",X"77",X"47",X"23",X"7E",
		X"90",X"D0",X"7E",X"4F",X"E6",X"F0",X"C6",X"10",X"2B",X"ED",X"44",X"86",X"77",X"79",X"E6",X"0F",
		X"FE",X"0F",X"20",X"38",X"18",X"34",X"3A",X"10",X"88",X"21",X"2A",X"88",X"0F",X"CB",X"16",X"7E",
		X"E6",X"07",X"FE",X"01",X"C0",X"EB",X"CD",X"09",X"0F",X"21",X"24",X"88",X"34",X"EB",X"23",X"7E",
		X"C6",X"10",X"77",X"47",X"23",X"7E",X"90",X"D0",X"7E",X"4F",X"E6",X"F0",X"C6",X"10",X"2B",X"ED",
		X"44",X"86",X"77",X"79",X"E6",X"0F",X"FE",X"0F",X"20",X"02",X"3E",X"63",X"21",X"02",X"88",X"86",
		X"77",X"FE",X"63",X"38",X"02",X"36",X"63",X"11",X"01",X"07",X"FF",X"C9",X"3A",X"24",X"88",X"A7",
		X"C8",X"21",X"25",X"88",X"7E",X"A7",X"20",X"07",X"36",X"30",X"3C",X"32",X"83",X"A1",X"C9",X"35",
		X"28",X"09",X"7E",X"FE",X"18",X"C0",X"AF",X"32",X"83",X"A1",X"C9",X"21",X"24",X"88",X"35",X"C9",
		X"3A",X"26",X"88",X"A7",X"C8",X"21",X"27",X"88",X"7E",X"A7",X"20",X"07",X"36",X"30",X"3C",X"32",
		X"84",X"A1",X"C9",X"35",X"28",X"09",X"7E",X"FE",X"18",X"C0",X"AF",X"32",X"84",X"A1",X"C9",X"21",
		X"26",X"88",X"35",X"C9",X"CD",X"78",X"5E",X"CD",X"6A",X"5F",X"CD",X"2F",X"60",X"CD",X"68",X"63",
		X"CD",X"F7",X"5D",X"CD",X"06",X"5B",X"CD",X"4D",X"5D",X"CD",X"86",X"5B",X"CD",X"04",X"64",X"CD",
		X"0B",X"5D",X"CD",X"2C",X"5B",X"C9",X"3A",X"07",X"89",X"FE",X"05",X"C0",X"FD",X"21",X"15",X"53",
		X"FD",X"55",X"FD",X"5C",X"AF",X"6F",X"67",X"06",X"06",X"1A",X"85",X"30",X"01",X"24",X"6F",X"13",
		X"10",X"F7",X"84",X"C6",X"7F",X"C8",X"26",X"88",X"2E",X"1E",X"34",X"C9",X"3A",X"75",X"8D",X"A7",
		X"C8",X"3A",X"79",X"8D",X"A7",X"C0",X"3A",X"77",X"8D",X"A7",X"20",X"1B",X"21",X"E4",X"8A",X"11",
		X"18",X"00",X"06",X"06",X"0E",X"13",X"3A",X"07",X"89",X"CB",X"47",X"28",X"02",X"0E",X"0B",X"7E",
		X"B9",X"28",X"04",X"19",X"10",X"F9",X"C9",X"DD",X"21",X"E0",X"8A",X"11",X"18",X"00",X"06",X"06",
		X"D9",X"CD",X"71",X"5B",X"D9",X"DD",X"19",X"10",X"F7",X"AF",X"32",X"75",X"8D",X"32",X"20",X"8F",
		X"C9",X"DD",X"7E",X"02",X"FE",X"05",X"C0",X"DD",X"CB",X"07",X"56",X"C8",X"DD",X"7E",X"06",X"FE",
		X"11",X"D0",X"CD",X"6C",X"3A",X"C9",X"DD",X"21",X"E0",X"8A",X"11",X"18",X"00",X"06",X"06",X"D9",
		X"CD",X"99",X"5B",X"D9",X"DD",X"19",X"10",X"F7",X"C9",X"DD",X"CB",X"0B",X"46",X"20",X"06",X"3A",
		X"07",X"89",X"CB",X"47",X"C0",X"DD",X"CB",X"00",X"46",X"C8",X"DD",X"CB",X"16",X"46",X"C8",X"DD",
		X"7E",X"02",X"FE",X"05",X"C0",X"21",X"48",X"88",X"FD",X"21",X"90",X"8C",X"06",X"02",X"FD",X"CB",
		X"00",X"46",X"CA",X"46",X"5C",X"FD",X"CB",X"00",X"4E",X"20",X"7B",X"1E",X"10",X"3A",X"1F",X"88",
		X"A7",X"20",X"02",X"1E",X"08",X"DD",X"7E",X"06",X"DD",X"4E",X"05",X"CB",X"01",X"17",X"CB",X"01",
		X"17",X"CB",X"01",X"17",X"83",X"FD",X"96",X"06",X"30",X"02",X"ED",X"44",X"FE",X"10",X"30",X"56",
		X"2C",X"2C",X"1E",X"16",X"3A",X"07",X"89",X"CB",X"47",X"20",X"02",X"1E",X"12",X"DD",X"7E",X"04",
		X"DD",X"4E",X"03",X"CB",X"01",X"17",X"CB",X"01",X"17",X"CB",X"01",X"17",X"93",X"FD",X"96",X"04",
		X"30",X"02",X"ED",X"44",X"FE",X"09",X"30",X"30",X"11",X"80",X"5C",X"DD",X"CB",X"07",X"4E",X"28",
		X"03",X"11",X"89",X"5C",X"CD",X"1E",X"38",X"DD",X"36",X"12",X"10",X"DD",X"36",X"16",X"02",X"FD",
		X"21",X"70",X"8B",X"11",X"18",X"00",X"06",X"05",X"DD",X"7E",X"14",X"FD",X"BE",X"14",X"28",X"14",
		X"FD",X"19",X"10",X"F4",X"F1",X"C9",X"2C",X"2C",X"2C",X"2C",X"11",X"18",X"00",X"FD",X"19",X"05",
		X"C2",X"BE",X"5B",X"C9",X"21",X"92",X"5C",X"DD",X"7E",X"07",X"E6",X"F0",X"0F",X"0F",X"0F",X"0F",
		X"CD",X"45",X"0C",X"FD",X"CB",X"0B",X"46",X"28",X"03",X"11",X"F9",X"5C",X"FD",X"36",X"16",X"02",
		X"CD",X"75",X"5C",X"F1",X"C9",X"FD",X"73",X"0C",X"FD",X"72",X"0D",X"FD",X"36",X"0E",X"00",X"C9",
		X"80",X"01",X"10",X"40",X"29",X"F0",X"FF",X"83",X"5C",X"84",X"01",X"10",X"44",X"29",X"F0",X"FF",
		X"8C",X"5C",X"A8",X"5C",X"B1",X"5C",X"BA",X"5C",X"C3",X"5C",X"CC",X"5C",X"D5",X"5C",X"DE",X"5C",
		X"DE",X"5C",X"DE",X"5C",X"E7",X"5C",X"F0",X"5C",X"40",X"20",X"10",X"40",X"22",X"F0",X"FF",X"AB",
		X"5C",X"41",X"20",X"10",X"41",X"22",X"F0",X"FF",X"B4",X"5C",X"44",X"20",X"10",X"44",X"22",X"F0",
		X"FF",X"BD",X"5C",X"49",X"20",X"10",X"49",X"22",X"F0",X"FF",X"C6",X"5C",X"4A",X"20",X"10",X"4A",
		X"22",X"F0",X"FF",X"CF",X"5C",X"41",X"20",X"10",X"41",X"22",X"F0",X"FF",X"D8",X"5C",X"44",X"20",
		X"10",X"44",X"22",X"F0",X"FF",X"E1",X"5C",X"4E",X"20",X"10",X"4E",X"22",X"F0",X"FF",X"EA",X"5C",
		X"4F",X"20",X"10",X"4F",X"22",X"F0",X"FF",X"F3",X"5C",X"44",X"20",X"10",X"44",X"A1",X"08",X"4B",
		X"A1",X"08",X"4C",X"A1",X"08",X"4F",X"A1",X"08",X"FF",X"FC",X"5C",X"DD",X"21",X"E0",X"8A",X"11",
		X"18",X"00",X"06",X"06",X"D9",X"CD",X"1E",X"5D",X"D9",X"DD",X"19",X"10",X"F7",X"C9",X"DD",X"CB",
		X"0B",X"46",X"20",X"06",X"3A",X"07",X"89",X"CB",X"47",X"C0",X"DD",X"CB",X"00",X"46",X"C8",X"DD",
		X"CB",X"16",X"4E",X"C8",X"DD",X"35",X"12",X"C0",X"DD",X"7E",X"13",X"E6",X"03",X"28",X"09",X"3D",
		X"DD",X"77",X"13",X"DD",X"36",X"16",X"01",X"C9",X"DD",X"36",X"16",X"00",X"C9",X"DD",X"21",X"9C",
		X"88",X"FD",X"21",X"7C",X"88",X"21",X"E8",X"8B",X"06",X"03",X"CD",X"68",X"5D",X"11",X"04",X"00",
		X"FD",X"19",X"1E",X"18",X"19",X"10",X"F3",X"C9",X"7E",X"A7",X"C8",X"FE",X"05",X"C8",X"1E",X"FC",
		X"16",X"00",X"3A",X"1F",X"88",X"A7",X"20",X"04",X"1E",X"05",X"16",X"10",X"DD",X"7E",X"00",X"83",
		X"5F",X"DD",X"7E",X"02",X"82",X"57",X"FD",X"7E",X"00",X"93",X"30",X"02",X"ED",X"44",X"FE",X"04",
		X"D0",X"FD",X"7E",X"02",X"C6",X"08",X"92",X"30",X"02",X"ED",X"44",X"FE",X"09",X"D8",X"FE",X"0F",
		X"D0",X"E5",X"DD",X"E1",X"DD",X"36",X"00",X"00",X"DD",X"36",X"01",X"01",X"DD",X"36",X"02",X"0C",
		X"DD",X"36",X"07",X"01",X"21",X"C2",X"5D",X"DD",X"74",X"13",X"DD",X"75",X"12",X"CD",X"2B",X"0F",
		X"F1",X"C9",X"60",X"20",X"60",X"20",X"40",X"20",X"40",X"40",X"40",X"40",X"40",X"40",X"20",X"40",
		X"20",X"40",X"20",X"40",X"20",X"60",X"20",X"60",X"20",X"40",X"20",X"60",X"20",X"60",X"20",X"60",
		X"20",X"60",X"20",X"60",X"20",X"60",X"20",X"60",X"20",X"60",X"20",X"60",X"10",X"60",X"10",X"60",
		X"10",X"60",X"10",X"60",X"EE",X"0C",X"60",X"3A",X"32",X"8D",X"A7",X"C0",X"3A",X"08",X"8F",X"21",
		X"24",X"8F",X"B6",X"C0",X"DD",X"21",X"40",X"88",X"FD",X"21",X"7C",X"88",X"21",X"E8",X"8B",X"06",
		X"03",X"CD",X"1F",X"5E",X"11",X"04",X"00",X"FD",X"19",X"1E",X"18",X"19",X"10",X"F3",X"C9",X"7E",
		X"A7",X"C8",X"FE",X"05",X"C8",X"1E",X"09",X"16",X"00",X"3A",X"1F",X"88",X"A7",X"20",X"04",X"1E",
		X"F7",X"16",X"10",X"DD",X"7E",X"00",X"83",X"5F",X"DD",X"7E",X"02",X"82",X"57",X"FD",X"7E",X"00",
		X"93",X"30",X"02",X"ED",X"44",X"FE",X"02",X"D0",X"FD",X"7E",X"02",X"C6",X"08",X"92",X"30",X"02",
		X"ED",X"44",X"FE",X"09",X"D0",X"3E",X"01",X"32",X"32",X"8D",X"E5",X"DD",X"E1",X"11",X"B4",X"40",
		X"CD",X"1E",X"38",X"DD",X"36",X"11",X"0A",X"DD",X"36",X"00",X"00",X"DD",X"36",X"01",X"01",X"DD",
		X"36",X"02",X"02",X"CD",X"15",X"0F",X"F1",X"C9",X"3A",X"07",X"89",X"E6",X"01",X"C8",X"FD",X"21",
		X"48",X"88",X"06",X"02",X"11",X"04",X"00",X"AF",X"ED",X"47",X"D9",X"CD",X"98",X"5E",X"D9",X"FD",
		X"19",X"3E",X"01",X"ED",X"47",X"10",X"F3",X"C9",X"ED",X"57",X"DD",X"21",X"90",X"8C",X"A7",X"28",
		X"04",X"DD",X"21",X"A8",X"8C",X"DD",X"CB",X"00",X"46",X"C8",X"DD",X"22",X"65",X"8D",X"DD",X"CB",
		X"00",X"4E",X"DD",X"21",X"88",X"88",X"06",X"04",X"21",X"30",X"8C",X"20",X"54",X"7E",X"A7",X"28",
		X"45",X"2C",X"2C",X"7E",X"2D",X"2D",X"FE",X"04",X"30",X"3C",X"CD",X"53",X"5F",X"30",X"37",X"57",
		X"FD",X"7E",X"00",X"93",X"30",X"02",X"ED",X"44",X"FE",X"0A",X"30",X"2A",X"FD",X"7E",X"02",X"C6",
		X"08",X"92",X"30",X"02",X"ED",X"44",X"FE",X"09",X"30",X"1C",X"AF",X"77",X"23",X"36",X"01",X"23",
		X"36",X"08",X"DD",X"2A",X"65",X"8D",X"DD",X"CB",X"07",X"46",X"20",X"06",X"2A",X"65",X"8D",X"06",
		X"17",X"D7",X"CD",X"F1",X"0E",X"C9",X"11",X"04",X"00",X"DD",X"19",X"1E",X"18",X"19",X"10",X"AD",
		X"C9",X"7E",X"A7",X"28",X"32",X"FE",X"03",X"28",X"2E",X"CD",X"53",X"5F",X"30",X"29",X"57",X"FD",
		X"7E",X"00",X"93",X"30",X"02",X"ED",X"44",X"FE",X"07",X"30",X"1C",X"FD",X"7E",X"02",X"C6",X"08",
		X"92",X"30",X"02",X"ED",X"44",X"FE",X"06",X"30",X"0E",X"36",X"03",X"21",X"19",X"8D",X"ED",X"57",
		X"28",X"01",X"2C",X"36",X"01",X"18",X"BB",X"11",X"04",X"00",X"DD",X"19",X"11",X"18",X"00",X"19",
		X"10",X"BF",X"C9",X"1E",X"06",X"3A",X"1F",X"88",X"A7",X"20",X"02",X"1E",X"FE",X"DD",X"7E",X"00",
		X"83",X"5F",X"DD",X"7E",X"02",X"C6",X"08",X"FE",X"E0",X"C9",X"FD",X"21",X"48",X"88",X"06",X"02",
		X"11",X"04",X"00",X"AF",X"ED",X"47",X"D9",X"CD",X"83",X"5F",X"D9",X"FD",X"19",X"78",X"ED",X"47",
		X"10",X"F4",X"C9",X"DD",X"21",X"90",X"8C",X"ED",X"57",X"A7",X"28",X"04",X"DD",X"21",X"A8",X"8C",
		X"DD",X"7E",X"00",X"A7",X"C8",X"32",X"44",X"8D",X"4F",X"DD",X"21",X"50",X"88",X"06",X"06",X"21",
		X"E0",X"8A",X"7E",X"A7",X"28",X"72",X"2C",X"2C",X"7E",X"2D",X"2D",X"FE",X"05",X"20",X"69",X"1E",
		X"06",X"3A",X"1F",X"88",X"A7",X"20",X"02",X"1E",X"FB",X"DD",X"7E",X"00",X"83",X"5F",X"DD",X"7E",
		X"02",X"C6",X"08",X"57",X"FD",X"7E",X"00",X"93",X"30",X"02",X"ED",X"44",X"5F",X"79",X"FE",X"03",
		X"7B",X"20",X"06",X"FE",X"10",X"30",X"41",X"18",X"04",X"FE",X"08",X"30",X"3B",X"FD",X"7E",X"02",
		X"C6",X"08",X"92",X"30",X"02",X"ED",X"44",X"5F",X"79",X"FE",X"03",X"7B",X"20",X"06",X"FE",X"12",
		X"30",X"26",X"18",X"04",X"FE",X"08",X"30",X"20",X"79",X"FE",X"03",X"28",X"28",X"FD",X"E5",X"E1",
		X"7D",X"21",X"91",X"8C",X"FE",X"48",X"28",X"03",X"21",X"A9",X"8C",X"36",X"01",X"11",X"06",X"00",
		X"19",X"36",X"01",X"CD",X"01",X"0F",X"F1",X"C9",X"11",X"04",X"00",X"DD",X"19",X"1E",X"18",X"19",
		X"05",X"C2",X"A2",X"5F",X"C9",X"E5",X"FD",X"E1",X"21",X"45",X"8D",X"34",X"C3",X"3D",X"61",X"FD",
		X"21",X"48",X"88",X"06",X"02",X"AF",X"ED",X"47",X"11",X"04",X"00",X"D9",X"CD",X"48",X"60",X"D9",
		X"FD",X"19",X"78",X"ED",X"47",X"10",X"F4",X"C9",X"DD",X"21",X"90",X"8C",X"ED",X"57",X"A7",X"28",
		X"04",X"DD",X"21",X"A8",X"8C",X"DD",X"7E",X"00",X"A7",X"C8",X"FE",X"03",X"C8",X"32",X"44",X"8D",
		X"DD",X"21",X"68",X"88",X"06",X"05",X"21",X"70",X"8B",X"7E",X"A7",X"CA",X"F2",X"60",X"2C",X"2C",
		X"7E",X"2D",X"2D",X"FE",X"05",X"C2",X"F2",X"60",X"3A",X"07",X"89",X"CB",X"47",X"C2",X"B4",X"61",
		X"1E",X"06",X"3A",X"1F",X"88",X"A7",X"20",X"02",X"1E",X"FE",X"DD",X"7E",X"00",X"83",X"5F",X"DD",
		X"7E",X"02",X"C6",X"08",X"57",X"FD",X"7E",X"00",X"93",X"30",X"02",X"ED",X"44",X"FE",X"09",X"30",
		X"51",X"FD",X"7E",X"02",X"C6",X"08",X"92",X"30",X"02",X"ED",X"44",X"FE",X"08",X"30",X"43",X"11",
		X"14",X"00",X"19",X"FD",X"21",X"E0",X"8A",X"7E",X"0E",X"06",X"1E",X"18",X"FD",X"BE",X"14",X"28",
		X"07",X"FD",X"19",X"0D",X"20",X"F6",X"18",X"0D",X"FD",X"CB",X"16",X"4E",X"28",X"07",X"3A",X"44",
		X"8D",X"FE",X"03",X"20",X"2A",X"11",X"EC",X"FF",X"19",X"FD",X"21",X"1C",X"8D",X"ED",X"57",X"20",
		X"02",X"FD",X"2B",X"FD",X"36",X"00",X"01",X"11",X"04",X"04",X"CD",X"9F",X"61",X"11",X"FD",X"FF",
		X"18",X"2D",X"11",X"04",X"00",X"DD",X"19",X"1E",X"18",X"19",X"05",X"C2",X"69",X"60",X"C9",X"DD",
		X"21",X"90",X"8C",X"ED",X"57",X"28",X"04",X"DD",X"21",X"A8",X"8C",X"DD",X"36",X"01",X"01",X"DD",
		X"36",X"07",X"01",X"CD",X"01",X"0F",X"F1",X"C9",X"3A",X"45",X"8D",X"3C",X"32",X"45",X"8D",X"19",
		X"7E",X"06",X"06",X"11",X"18",X"00",X"FD",X"21",X"E0",X"8A",X"FD",X"BE",X"14",X"28",X"0E",X"FD",
		X"19",X"10",X"F7",X"3A",X"44",X"8D",X"FE",X"03",X"C8",X"CD",X"F1",X"0E",X"C9",X"FD",X"CB",X"00",
		X"46",X"28",X"47",X"3A",X"07",X"89",X"E6",X"01",X"20",X"1C",X"3A",X"44",X"8D",X"FE",X"03",X"20",
		X"15",X"FD",X"7E",X"14",X"DD",X"21",X"70",X"8B",X"11",X"18",X"00",X"06",X"06",X"DD",X"BE",X"14",
		X"28",X"2E",X"DD",X"19",X"10",X"F7",X"AF",X"FD",X"77",X"00",X"FD",X"36",X"01",X"01",X"FD",X"36",
		X"02",X"08",X"FD",X"36",X"16",X"07",X"FD",X"36",X"17",X"05",X"FD",X"77",X"14",X"FD",X"77",X"13",
		X"3A",X"44",X"8D",X"FE",X"03",X"20",X"13",X"CD",X"FD",X"0E",X"AF",X"32",X"44",X"8D",X"F1",X"C9",
		X"DD",X"36",X"08",X"01",X"DD",X"36",X"0A",X"D0",X"18",X"CC",X"CD",X"F1",X"0E",X"18",X"EB",X"36",
		X"00",X"23",X"36",X"01",X"23",X"36",X"08",X"01",X"10",X"00",X"09",X"36",X"FF",X"0E",X"04",X"09",
		X"73",X"23",X"72",X"C9",X"E5",X"FD",X"E5",X"C5",X"7D",X"C6",X"14",X"6F",X"7E",X"FD",X"21",X"E0",
		X"8A",X"01",X"18",X"00",X"2E",X"05",X"FD",X"BE",X"14",X"28",X"0C",X"FD",X"09",X"2D",X"20",X"F6",
		X"C1",X"FD",X"E1",X"E1",X"C3",X"80",X"60",X"FD",X"7E",X"0B",X"A7",X"20",X"F3",X"FD",X"7E",X"16",
		X"C1",X"FD",X"E1",X"E1",X"E6",X"F0",X"CA",X"80",X"60",X"FE",X"40",X"28",X"0F",X"FE",X"50",X"CA",
		X"87",X"62",X"FE",X"F0",X"CA",X"0F",X"63",X"FE",X"D0",X"CA",X"87",X"62",X"1E",X"06",X"3A",X"1F",
		X"88",X"A7",X"20",X"02",X"1E",X"FE",X"DD",X"7E",X"00",X"83",X"5F",X"DD",X"7E",X"02",X"C6",X"08",
		X"57",X"FD",X"7E",X"00",X"93",X"30",X"02",X"ED",X"44",X"FE",X"09",X"D2",X"F2",X"60",X"FD",X"7E",
		X"02",X"C6",X"08",X"92",X"30",X"02",X"ED",X"44",X"FE",X"08",X"D2",X"F2",X"60",X"E5",X"DD",X"E1",
		X"11",X"43",X"63",X"CD",X"1E",X"38",X"21",X"58",X"63",X"3A",X"07",X"89",X"E6",X"07",X"1F",X"E7",
		X"6F",X"DD",X"7E",X"0A",X"85",X"DD",X"77",X"0A",X"FD",X"21",X"E0",X"8A",X"DD",X"7E",X"14",X"0E",
		X"06",X"11",X"18",X"00",X"FD",X"BE",X"14",X"28",X"05",X"FD",X"19",X"0D",X"20",X"F6",X"21",X"58",
		X"63",X"3A",X"07",X"89",X"E6",X"07",X"1F",X"E7",X"6F",X"FD",X"7E",X"0A",X"85",X"FD",X"77",X"0A",
		X"FD",X"CB",X"16",X"E6",X"21",X"90",X"8C",X"ED",X"57",X"28",X"03",X"21",X"A8",X"8C",X"06",X"18",
		X"AF",X"D7",X"CD",X"F1",X"0E",X"F1",X"C9",X"4F",X"1E",X"06",X"3A",X"1F",X"88",X"A7",X"20",X"02",
		X"1E",X"FE",X"DD",X"7E",X"00",X"83",X"5F",X"DD",X"7E",X"02",X"C6",X"08",X"57",X"FD",X"7E",X"00",
		X"93",X"30",X"02",X"ED",X"44",X"FE",X"06",X"D2",X"F2",X"60",X"FD",X"7E",X"02",X"C6",X"08",X"92",
		X"30",X"02",X"ED",X"44",X"FE",X"07",X"D2",X"F2",X"60",X"79",X"FE",X"50",X"CA",X"D9",X"60",X"E5",
		X"DD",X"E1",X"11",X"49",X"63",X"CD",X"1E",X"38",X"21",X"60",X"63",X"3A",X"07",X"89",X"E6",X"07",
		X"1F",X"E7",X"6F",X"DD",X"7E",X"0A",X"85",X"DD",X"77",X"0A",X"FD",X"21",X"E0",X"8A",X"DD",X"7E",
		X"14",X"0E",X"06",X"11",X"18",X"00",X"FD",X"BE",X"14",X"28",X"05",X"FD",X"19",X"0D",X"20",X"F6",
		X"21",X"60",X"63",X"3A",X"07",X"89",X"E6",X"07",X"1F",X"E7",X"6F",X"FD",X"7E",X"0A",X"85",X"FD",
		X"77",X"0A",X"FD",X"CB",X"16",X"EE",X"11",X"4F",X"63",X"CD",X"75",X"5C",X"C3",X"74",X"62",X"1E",
		X"06",X"3A",X"1F",X"88",X"A7",X"20",X"02",X"1E",X"FE",X"DD",X"7E",X"00",X"83",X"5F",X"DD",X"7E",
		X"02",X"C6",X"08",X"57",X"FD",X"7E",X"00",X"93",X"30",X"02",X"ED",X"44",X"FE",X"05",X"D2",X"F2",
		X"60",X"FD",X"7E",X"02",X"C6",X"08",X"92",X"30",X"02",X"ED",X"44",X"FE",X"05",X"D2",X"F2",X"60",
		X"C3",X"D9",X"60",X"41",X"23",X"F0",X"FF",X"43",X"63",X"4C",X"24",X"F0",X"FF",X"49",X"63",X"40",
		X"0B",X"0D",X"40",X"06",X"0D",X"FF",X"4F",X"63",X"08",X"09",X"0A",X"0B",X"0C",X"0D",X"0E",X"0E",
		X"06",X"07",X"08",X"09",X"0A",X"0B",X"0C",X"0C",X"FD",X"21",X"48",X"88",X"06",X"02",X"11",X"04",
		X"00",X"AF",X"ED",X"47",X"D9",X"CD",X"81",X"63",X"D9",X"FD",X"19",X"7B",X"ED",X"47",X"10",X"F4",
		X"C9",X"DD",X"21",X"7C",X"88",X"06",X"03",X"21",X"E8",X"8B",X"7E",X"A7",X"28",X"61",X"1E",X"05",
		X"3A",X"1F",X"88",X"A7",X"20",X"02",X"1E",X"FE",X"DD",X"7E",X"00",X"83",X"5F",X"DD",X"7E",X"02",
		X"C6",X"08",X"57",X"FD",X"7E",X"00",X"93",X"30",X"02",X"ED",X"44",X"FE",X"06",X"30",X"40",X"FD",
		X"7E",X"02",X"C6",X"08",X"92",X"30",X"02",X"ED",X"44",X"FE",X"06",X"30",X"32",X"E5",X"DD",X"E1",
		X"DD",X"36",X"00",X"00",X"DD",X"36",X"01",X"01",X"DD",X"36",X"02",X"02",X"DD",X"36",X"11",X"28",
		X"11",X"0F",X"00",X"21",X"1B",X"8D",X"ED",X"57",X"A7",X"28",X"03",X"21",X"1C",X"8D",X"36",X"01",
		X"11",X"FB",X"63",X"CD",X"1E",X"38",X"CD",X"F9",X"0E",X"11",X"15",X"03",X"FF",X"F1",X"C9",X"11",
		X"04",X"00",X"DD",X"19",X"11",X"18",X"00",X"19",X"10",X"90",X"C9",X"4F",X"34",X"06",X"4F",X"33",
		X"06",X"42",X"37",X"28",X"3A",X"50",X"8F",X"A7",X"20",X"06",X"3A",X"07",X"89",X"E6",X"01",X"C0",
		X"FD",X"21",X"48",X"88",X"06",X"02",X"11",X"04",X"00",X"AF",X"ED",X"47",X"D9",X"CD",X"35",X"64",
		X"D9",X"FD",X"19",X"7B",X"ED",X"47",X"10",X"F4",X"C9",X"11",X"04",X"00",X"DD",X"19",X"11",X"18",
		X"00",X"19",X"10",X"17",X"C9",X"DD",X"21",X"8C",X"88",X"21",X"48",X"8C",X"3A",X"50",X"8F",X"A7",
		X"28",X"07",X"DD",X"21",X"7C",X"88",X"21",X"E8",X"8B",X"06",X"03",X"7E",X"A7",X"28",X"DA",X"1E",
		X"05",X"3A",X"1F",X"88",X"A7",X"20",X"02",X"1E",X"FE",X"DD",X"7E",X"00",X"83",X"5F",X"DD",X"7E",
		X"02",X"C6",X"08",X"57",X"FD",X"7E",X"00",X"93",X"30",X"02",X"ED",X"44",X"FE",X"07",X"30",X"B9",
		X"FD",X"7E",X"02",X"C6",X"08",X"92",X"30",X"02",X"ED",X"44",X"FE",X"07",X"30",X"AB",X"E5",X"DD",
		X"E1",X"DD",X"36",X"00",X"00",X"DD",X"36",X"01",X"01",X"DD",X"36",X"02",X"02",X"DD",X"36",X"11",
		X"20",X"11",X"0F",X"00",X"21",X"1B",X"8D",X"ED",X"57",X"A7",X"28",X"03",X"21",X"1C",X"8D",X"36",
		X"01",X"11",X"DF",X"64",X"CD",X"1E",X"38",X"CD",X"F5",X"0E",X"3A",X"50",X"8F",X"A7",X"20",X"04",
		X"11",X"15",X"03",X"FF",X"21",X"52",X"8F",X"34",X"11",X"C2",X"0B",X"21",X"D0",X"64",X"1A",X"96",
		X"20",X"08",X"1B",X"23",X"7E",X"3D",X"28",X"06",X"18",X"F4",X"21",X"F9",X"8D",X"34",X"F1",X"C9",
		X"51",X"3A",X"3B",X"20",X"3D",X"88",X"05",X"3A",X"41",X"20",X"A7",X"88",X"06",X"3A",X"01",X"42",
		X"37",X"28",X"CD",X"13",X"6B",X"DD",X"21",X"78",X"8C",X"CD",X"FB",X"64",X"DD",X"21",X"E0",X"8A",
		X"FD",X"21",X"78",X"8C",X"CD",X"C5",X"66",X"CD",X"22",X"68",X"C9",X"DD",X"7E",X"02",X"EF",X"05",
		X"65",X"66",X"65",X"66",X"66",X"21",X"29",X"89",X"36",X"1C",X"11",X"E8",X"FF",X"06",X"03",X"2E",
		X"2B",X"36",X"08",X"D9",X"CD",X"23",X"65",X"D9",X"DD",X"34",X"02",X"DD",X"19",X"10",X"F4",X"CD",
		X"88",X"0F",X"C9",X"DD",X"7E",X"00",X"DD",X"B6",X"01",X"0F",X"D8",X"3A",X"F0",X"8E",X"A7",X"C0",
		X"DD",X"36",X"00",X"01",X"DD",X"77",X"03",X"DD",X"77",X"05",X"DD",X"36",X"04",X"15",X"3A",X"29",
		X"89",X"DD",X"77",X"06",X"D6",X"02",X"32",X"29",X"89",X"DD",X"36",X"0F",X"03",X"DD",X"36",X"10",
		X"C0",X"DD",X"36",X"08",X"30",X"DD",X"36",X"09",X"F0",X"11",X"11",X"06",X"FF",X"3A",X"07",X"89",
		X"A7",X"C0",X"1E",X"07",X"FF",X"C9",X"21",X"2F",X"89",X"7E",X"A7",X"28",X"02",X"35",X"C9",X"2E",
		X"2C",X"34",X"CB",X"46",X"2E",X"2F",X"20",X"1E",X"36",X"06",X"DD",X"7E",X"03",X"DD",X"86",X"08",
		X"30",X"09",X"DD",X"34",X"04",X"DD",X"34",X"EC",X"DD",X"34",X"D4",X"DD",X"77",X"03",X"DD",X"77",
		X"EB",X"DD",X"77",X"D3",X"18",X"54",X"36",X"0C",X"DD",X"7E",X"03",X"DD",X"96",X"08",X"30",X"09",
		X"DD",X"35",X"04",X"DD",X"35",X"EC",X"DD",X"35",X"D4",X"DD",X"77",X"03",X"DD",X"77",X"EB",X"DD",
		X"77",X"D3",X"DD",X"7E",X"05",X"DD",X"96",X"09",X"DD",X"77",X"05",X"DD",X"77",X"ED",X"DD",X"77",
		X"D5",X"30",X"12",X"DD",X"7E",X"06",X"D6",X"01",X"DD",X"77",X"06",X"D6",X"02",X"DD",X"77",X"EE",
		X"D6",X"02",X"DD",X"77",X"D6",X"2E",X"2C",X"CB",X"46",X"21",X"BF",X"66",X"28",X"03",X"21",X"C2",
		X"66",X"11",X"E8",X"FF",X"06",X"03",X"CD",X"14",X"25",X"C9",X"DD",X"21",X"78",X"8C",X"DD",X"7E",
		X"06",X"FE",X"0C",X"D0",X"3E",X"40",X"DD",X"77",X"10",X"DD",X"77",X"F8",X"DD",X"77",X"E0",X"3E",
		X"18",X"DD",X"77",X"09",X"DD",X"77",X"F1",X"DD",X"77",X"D9",X"3E",X"02",X"DD",X"77",X"02",X"DD",
		X"77",X"EA",X"DD",X"77",X"D2",X"32",X"30",X"89",X"32",X"2E",X"89",X"FD",X"21",X"BC",X"82",X"11",
		X"00",X"00",X"06",X"0A",X"FD",X"7E",X"00",X"FD",X"BE",X"E0",X"C2",X"84",X"52",X"83",X"5F",X"30",
		X"01",X"14",X"FD",X"7D",X"D6",X"20",X"FD",X"6F",X"30",X"02",X"FD",X"25",X"10",X"E6",X"06",X"0A",
		X"3E",X"04",X"FD",X"84",X"FD",X"67",X"EB",X"FD",X"5D",X"FD",X"54",X"EB",X"7E",X"83",X"30",X"01",
		X"14",X"5F",X"7D",X"C6",X"20",X"30",X"01",X"24",X"6F",X"10",X"F1",X"7B",X"FE",X"2A",X"C2",X"14",
		X"60",X"15",X"C2",X"05",X"20",X"C9",X"11",X"E8",X"FF",X"06",X"03",X"D9",X"CD",X"7C",X"66",X"D9",
		X"DD",X"19",X"10",X"F7",X"DD",X"21",X"78",X"8C",X"CD",X"A1",X"66",X"C9",X"DD",X"7E",X"01",X"A7",
		X"C0",X"DD",X"7E",X"05",X"DD",X"86",X"09",X"30",X"03",X"DD",X"34",X"06",X"DD",X"77",X"05",X"DD",
		X"7E",X"06",X"FE",X"1D",X"D8",X"DD",X"36",X"01",X"02",X"AF",X"DD",X"77",X"04",X"DD",X"77",X"06",
		X"C9",X"21",X"2B",X"89",X"35",X"7E",X"A7",X"C0",X"36",X"08",X"23",X"34",X"CB",X"46",X"21",X"BF",
		X"66",X"28",X"03",X"21",X"C2",X"66",X"11",X"E8",X"FF",X"06",X"03",X"CD",X"14",X"25",X"C9",X"03",
		X"03",X"03",X"09",X"09",X"09",X"11",X"18",X"00",X"06",X"03",X"D9",X"CD",X"F1",X"66",X"D9",X"DD",
		X"19",X"10",X"F7",X"3A",X"E2",X"8A",X"A7",X"C8",X"21",X"2D",X"89",X"7E",X"A7",X"28",X"02",X"35",
		X"C9",X"36",X"10",X"23",X"23",X"34",X"CB",X"46",X"11",X"12",X"06",X"20",X"02",X"1E",X"92",X"FF",
		X"C9",X"DD",X"7E",X"02",X"EF",X"FD",X"66",X"2A",X"67",X"A0",X"67",X"DF",X"67",X"3A",X"30",X"89",
		X"A7",X"C8",X"21",X"2E",X"89",X"7E",X"A7",X"28",X"02",X"35",X"C9",X"36",X"12",X"DD",X"34",X"02",
		X"AF",X"DD",X"77",X"03",X"DD",X"77",X"05",X"DD",X"36",X"04",X"15",X"DD",X"36",X"06",X"02",X"11",
		X"29",X"38",X"CD",X"1E",X"38",X"DD",X"36",X"09",X"2C",X"C9",X"CD",X"06",X"40",X"DD",X"7E",X"05",
		X"DD",X"86",X"09",X"30",X"03",X"DD",X"34",X"06",X"DD",X"77",X"05",X"DD",X"7E",X"06",X"FE",X"18",
		X"30",X"50",X"FD",X"21",X"48",X"8C",X"11",X"18",X"00",X"06",X"03",X"FD",X"7E",X"01",X"A7",X"20",
		X"08",X"DD",X"7E",X"06",X"FD",X"BE",X"06",X"28",X"05",X"FD",X"19",X"10",X"EE",X"C9",X"21",X"03",
		X"89",X"34",X"FD",X"36",X"01",X"02",X"DD",X"7E",X"03",X"D6",X"80",X"30",X"03",X"FD",X"35",X"04",
		X"FD",X"77",X"03",X"DD",X"7E",X"05",X"C6",X"40",X"30",X"03",X"FD",X"35",X"06",X"FD",X"77",X"05",
		X"FD",X"36",X"0F",X"C0",X"FD",X"E5",X"E1",X"DD",X"75",X"07",X"DD",X"74",X"08",X"3E",X"20",X"32",
		X"29",X"89",X"DD",X"34",X"02",X"DD",X"36",X"09",X"18",X"11",X"38",X"38",X"CD",X"1E",X"38",X"C9",
		X"21",X"29",X"89",X"7E",X"A7",X"28",X"02",X"35",X"C9",X"CD",X"06",X"40",X"DD",X"6E",X"07",X"DD",
		X"66",X"08",X"7C",X"A7",X"28",X"11",X"E5",X"FD",X"E1",X"FD",X"7E",X"05",X"DD",X"96",X"09",X"30",
		X"03",X"FD",X"35",X"06",X"FD",X"77",X"05",X"DD",X"7E",X"05",X"DD",X"96",X"09",X"30",X"03",X"DD",
		X"35",X"06",X"DD",X"77",X"05",X"DD",X"7E",X"06",X"FE",X"00",X"C0",X"DD",X"34",X"02",X"C9",X"21",
		X"BC",X"82",X"11",X"E0",X"FF",X"01",X"00",X"0A",X"7E",X"81",X"4F",X"19",X"10",X"FA",X"3E",X"5A",
		X"B9",X"20",X"AD",X"3E",X"01",X"32",X"04",X"89",X"32",X"08",X"88",X"32",X"0A",X"88",X"AF",X"21",
		X"28",X"89",X"06",X"09",X"D7",X"21",X"80",X"8A",X"77",X"11",X"81",X"8A",X"01",X"40",X"02",X"ED",
		X"B0",X"3E",X"10",X"21",X"42",X"84",X"0E",X"1D",X"06",X"1D",X"D7",X"23",X"23",X"23",X"0D",X"20",
		X"F7",X"C9",X"3A",X"FA",X"8A",X"A7",X"C8",X"DD",X"21",X"E0",X"8A",X"11",X"48",X"00",X"DD",X"19",
		X"DD",X"7E",X"02",X"EF",X"3A",X"68",X"57",X"68",X"AC",X"68",X"DD",X"34",X"02",X"AF",X"DD",X"77",
		X"03",X"DD",X"77",X"05",X"DD",X"36",X"04",X"08",X"DD",X"36",X"06",X"1E",X"11",X"EF",X"68",X"CD",
		X"1E",X"38",X"DD",X"36",X"09",X"18",X"C9",X"CD",X"06",X"40",X"DD",X"7E",X"05",X"DD",X"96",X"09",
		X"30",X"03",X"DD",X"35",X"06",X"DD",X"77",X"05",X"DD",X"7E",X"06",X"FE",X"1B",X"D0",X"DD",X"34",
		X"02",X"21",X"BC",X"86",X"11",X"A3",X"68",X"01",X"00",X"08",X"1A",X"86",X"81",X"4F",X"13",X"7D",
		X"D6",X"20",X"30",X"01",X"25",X"6F",X"10",X"F2",X"06",X"08",X"7C",X"D6",X"04",X"67",X"7E",X"81",
		X"4F",X"7D",X"C6",X"20",X"30",X"01",X"24",X"10",X"F5",X"1A",X"81",X"C2",X"B3",X"08",X"11",X"13",
		X"06",X"FF",X"C9",X"16",X"10",X"05",X"01",X"02",X"0F",X"03",X"07",X"B8",X"21",X"55",X"8F",X"7E",
		X"A7",X"C0",X"34",X"21",X"02",X"84",X"11",X"00",X"00",X"7E",X"83",X"5F",X"30",X"01",X"14",X"2C",
		X"7D",X"E6",X"1F",X"FE",X"1F",X"20",X"F2",X"7D",X"C6",X"03",X"6F",X"30",X"EC",X"24",X"7C",X"FE",
		X"88",X"38",X"E6",X"21",X"EB",X"68",X"06",X"04",X"7B",X"BE",X"28",X"06",X"23",X"10",X"FA",X"C3",
		X"D4",X"76",X"7A",X"23",X"BE",X"C8",X"10",X"FA",X"C3",X"29",X"38",X"43",X"95",X"89",X"87",X"40",
		X"15",X"08",X"40",X"1E",X"08",X"FF",X"EF",X"68",X"CD",X"05",X"69",X"CD",X"AD",X"69",X"CD",X"0F",
		X"6A",X"CD",X"7F",X"6A",X"C9",X"21",X"29",X"89",X"7E",X"A7",X"28",X"02",X"35",X"C9",X"2E",X"2D",
		X"7E",X"2E",X"03",X"BE",X"C8",X"FE",X"08",X"D0",X"DD",X"21",X"E0",X"8A",X"FD",X"21",X"A0",X"8B",
		X"11",X"18",X"00",X"06",X"08",X"D9",X"CD",X"31",X"69",X"D9",X"DD",X"19",X"FD",X"19",X"10",X"F5",
		X"C9",X"DD",X"7E",X"00",X"DD",X"B6",X"01",X"0F",X"D8",X"AF",X"DD",X"77",X"03",X"DD",X"77",X"05",
		X"3C",X"DD",X"77",X"00",X"FD",X"77",X"00",X"DD",X"36",X"04",X"15",X"DD",X"36",X"06",X"1E",X"FD",
		X"36",X"03",X"80",X"FD",X"36",X"05",X"A0",X"FD",X"36",X"04",X"14",X"FD",X"36",X"06",X"1E",X"FD",
		X"36",X"0F",X"03",X"FD",X"36",X"10",X"40",X"DD",X"36",X"09",X"24",X"FD",X"36",X"09",X"24",X"11",
		X"38",X"38",X"CD",X"1E",X"38",X"3E",X"10",X"32",X"29",X"89",X"3A",X"2D",X"89",X"A7",X"20",X"27",
		X"11",X"25",X"06",X"FF",X"1E",X"0A",X"FF",X"21",X"3B",X"86",X"3A",X"03",X"89",X"47",X"AF",X"C6",
		X"01",X"27",X"10",X"FB",X"5F",X"E6",X"F0",X"0F",X"0F",X"0F",X"0F",X"77",X"01",X"E0",X"FF",X"09",
		X"7B",X"E6",X"0F",X"77",X"CD",X"97",X"0F",X"21",X"2D",X"89",X"34",X"F1",X"C9",X"DD",X"21",X"E0",
		X"8A",X"FD",X"21",X"A0",X"8B",X"11",X"18",X"00",X"06",X"08",X"D9",X"CD",X"C6",X"69",X"D9",X"DD",
		X"19",X"FD",X"19",X"10",X"F5",X"C9",X"DD",X"7E",X"00",X"A7",X"C8",X"DD",X"7E",X"02",X"A7",X"C0",
		X"CD",X"06",X"40",X"FD",X"7E",X"05",X"FD",X"96",X"09",X"30",X"03",X"FD",X"35",X"06",X"FD",X"77",
		X"05",X"DD",X"7E",X"05",X"DD",X"96",X"09",X"30",X"03",X"DD",X"35",X"06",X"DD",X"77",X"05",X"DD",
		X"7E",X"06",X"FE",X"06",X"20",X"08",X"21",X"2B",X"89",X"7E",X"A7",X"C0",X"34",X"C9",X"FE",X"01",
		X"D0",X"AF",X"DD",X"E5",X"E1",X"06",X"18",X"D7",X"FD",X"E5",X"E1",X"06",X"18",X"D7",X"C9",X"21",
		X"2B",X"89",X"7E",X"A7",X"C8",X"23",X"7E",X"FE",X"06",X"C8",X"2E",X"2A",X"7E",X"A7",X"28",X"02",
		X"35",X"C9",X"DD",X"21",X"E0",X"8A",X"11",X"18",X"00",X"06",X"12",X"D9",X"CD",X"35",X"6A",X"D9",
		X"DD",X"19",X"10",X"F7",X"C9",X"DD",X"7E",X"00",X"DD",X"B6",X"01",X"0F",X"D8",X"AF",X"DD",X"77",
		X"03",X"DD",X"77",X"05",X"3C",X"DD",X"77",X"01",X"DD",X"77",X"02",X"DD",X"36",X"04",X"15",X"DD",
		X"36",X"06",X"1E",X"DD",X"36",X"09",X"28",X"21",X"2A",X"89",X"36",X"10",X"2E",X"2C",X"7E",X"34",
		X"FE",X"02",X"28",X"0E",X"30",X"11",X"A7",X"28",X"04",X"2E",X"2A",X"36",X"1C",X"11",X"D4",X"76",
		X"18",X"08",X"11",X"EF",X"68",X"18",X"03",X"11",X"0A",X"6B",X"CD",X"1E",X"38",X"F1",X"C9",X"3A",
		X"2B",X"89",X"A7",X"28",X"40",X"DD",X"21",X"E0",X"8A",X"11",X"18",X"00",X"06",X"12",X"D9",X"CD",
		X"98",X"6A",X"D9",X"DD",X"19",X"10",X"F7",X"C9",X"DD",X"7E",X"01",X"A7",X"C8",X"DD",X"7E",X"02",
		X"3D",X"E6",X"03",X"EF",X"A8",X"6A",X"DF",X"67",X"CD",X"06",X"40",X"DD",X"7E",X"05",X"DD",X"96",
		X"09",X"30",X"03",X"DD",X"35",X"06",X"DD",X"77",X"05",X"DD",X"7E",X"06",X"A7",X"C0",X"32",X"56",
		X"8F",X"DD",X"34",X"02",X"C9",X"3A",X"2D",X"89",X"FE",X"02",X"C0",X"3A",X"56",X"8F",X"A7",X"C0",
		X"3C",X"32",X"56",X"8F",X"21",X"50",X"84",X"11",X"00",X"00",X"7B",X"86",X"5F",X"30",X"01",X"14",
		X"2C",X"7D",X"E6",X"1F",X"FE",X"1B",X"20",X"03",X"2C",X"18",X"EF",X"FE",X"1F",X"20",X"EB",X"3E",
		X"12",X"85",X"6F",X"30",X"E5",X"24",X"7C",X"FE",X"88",X"38",X"DF",X"7B",X"FE",X"B8",X"28",X"03",
		X"C3",X"29",X"09",X"7A",X"FE",X"29",X"C2",X"29",X"38",X"C9",X"C0",X"03",X"08",X"C0",X"09",X"08",
		X"FF",X"0A",X"6B",X"21",X"06",X"8F",X"7E",X"A7",X"28",X"02",X"35",X"C9",X"36",X"0C",X"23",X"34",
		X"7E",X"E6",X"01",X"11",X"44",X"27",X"21",X"B4",X"84",X"28",X"03",X"11",X"48",X"27",X"D5",X"CD",
		X"25",X"33",X"11",X"A0",X"FF",X"19",X"D1",X"CD",X"25",X"33",X"C9",X"3A",X"06",X"88",X"A7",X"C0",
		X"3A",X"5F",X"8D",X"A7",X"C0",X"3A",X"07",X"89",X"E6",X"01",X"C0",X"21",X"5E",X"8D",X"7E",X"A7",
		X"C8",X"FE",X"01",X"28",X"02",X"35",X"C9",X"3E",X"11",X"32",X"0A",X"88",X"32",X"5F",X"8D",X"3E",
		X"FF",X"32",X"5E",X"8D",X"11",X"18",X"00",X"DD",X"21",X"E0",X"8A",X"FD",X"21",X"80",X"8D",X"06",
		X"0B",X"DD",X"7E",X"04",X"E6",X"1F",X"FE",X"06",X"38",X"1D",X"FE",X"1A",X"30",X"19",X"DD",X"E5",
		X"E1",X"FD",X"75",X"00",X"FD",X"74",X"01",X"DD",X"7E",X"06",X"FD",X"77",X"02",X"DD",X"36",X"06",
		X"00",X"FD",X"23",X"FD",X"23",X"FD",X"23",X"DD",X"19",X"10",X"D6",X"11",X"2B",X"06",X"FF",X"11",
		X"2C",X"06",X"FF",X"11",X"2D",X"06",X"FF",X"11",X"2E",X"06",X"FF",X"11",X"2F",X"06",X"FF",X"C3",
		X"EF",X"02",X"21",X"5E",X"8D",X"35",X"C0",X"FD",X"21",X"80",X"8D",X"11",X"03",X"00",X"06",X"0B",
		X"AF",X"FD",X"66",X"01",X"B4",X"28",X"09",X"FD",X"6E",X"00",X"FD",X"7E",X"02",X"19",X"19",X"77",
		X"FD",X"19",X"10",X"EC",X"3E",X"04",X"32",X"0A",X"88",X"11",X"AB",X"06",X"FF",X"11",X"AC",X"06",
		X"FF",X"11",X"AD",X"06",X"FF",X"11",X"AE",X"06",X"FF",X"11",X"AF",X"06",X"18",X"C0",X"3A",X"52",
		X"8D",X"A7",X"28",X"20",X"21",X"87",X"8A",X"3D",X"28",X"0D",X"CB",X"DE",X"CB",X"96",X"21",X"53",
		X"8D",X"35",X"C0",X"AF",X"2D",X"77",X"C9",X"CB",X"D6",X"CB",X"9E",X"21",X"53",X"8D",X"35",X"C0",
		X"AF",X"2D",X"77",X"C9",X"CD",X"18",X"6C",X"C9",X"DD",X"21",X"40",X"88",X"FD",X"21",X"7C",X"88",
		X"21",X"E8",X"8B",X"06",X"03",X"CD",X"3F",X"6C",X"11",X"04",X"00",X"FD",X"19",X"1E",X"18",X"19",
		X"10",X"F3",X"21",X"87",X"8A",X"CB",X"96",X"CB",X"9E",X"21",X"54",X"8D",X"36",X"00",X"C9",X"CB",
		X"46",X"C8",X"1E",X"10",X"16",X"00",X"DD",X"7E",X"00",X"83",X"5F",X"DD",X"7E",X"02",X"82",X"57",
		X"FD",X"7E",X"00",X"C6",X"20",X"93",X"30",X"02",X"ED",X"44",X"FE",X"18",X"D0",X"0E",X"00",X"FD",
		X"7E",X"02",X"C6",X"08",X"92",X"30",X"04",X"0E",X"FF",X"ED",X"44",X"FE",X"0E",X"D0",X"21",X"54",
		X"8D",X"36",X"01",X"DD",X"7E",X"02",X"21",X"87",X"8A",X"0C",X"20",X"13",X"FE",X"B6",X"38",X"1B",
		X"CB",X"D6",X"CB",X"9E",X"0E",X"01",X"21",X"52",X"8D",X"71",X"2C",X"36",X"18",X"F1",X"C9",X"FE",
		X"51",X"30",X"12",X"CB",X"DE",X"CB",X"96",X"0E",X"02",X"18",X"EB",X"FE",X"51",X"38",X"F4",X"CB",
		X"DE",X"CB",X"96",X"F1",X"C9",X"CB",X"D6",X"CB",X"9E",X"F1",X"C9",X"3A",X"06",X"88",X"A7",X"C0",
		X"3A",X"32",X"8D",X"A7",X"C0",X"3A",X"24",X"8F",X"A7",X"21",X"87",X"8A",X"28",X"03",X"AF",X"77",
		X"C9",X"CD",X"EE",X"6B",X"3A",X"54",X"8D",X"A7",X"C0",X"21",X"87",X"8A",X"3A",X"30",X"8F",X"FE",
		X"01",X"28",X"3A",X"3A",X"41",X"8F",X"A7",X"C2",X"4D",X"6D",X"21",X"42",X"88",X"DD",X"21",X"E0",
		X"8A",X"FD",X"21",X"52",X"88",X"06",X"06",X"DD",X"7E",X"00",X"A7",X"20",X"2A",X"11",X"18",X"00",
		X"DD",X"19",X"11",X"04",X"00",X"FD",X"19",X"10",X"EE",X"3A",X"41",X"8F",X"A7",X"C8",X"3A",X"42",
		X"88",X"4F",X"ED",X"5B",X"41",X"8F",X"21",X"87",X"8A",X"1A",X"B9",X"30",X"05",X"CB",X"D6",X"CB",
		X"9E",X"C9",X"CB",X"DE",X"CB",X"96",X"C9",X"FD",X"7E",X"00",X"FE",X"40",X"38",X"CF",X"FE",X"C0",
		X"30",X"CB",X"96",X"30",X"01",X"2F",X"4F",X"3A",X"40",X"8F",X"A7",X"28",X"04",X"B9",X"30",X"BD",
		X"79",X"32",X"40",X"8F",X"FD",X"E5",X"D1",X"7B",X"32",X"41",X"8F",X"7A",X"32",X"42",X"8F",X"DD",
		X"E5",X"D1",X"13",X"7B",X"32",X"43",X"8F",X"7A",X"32",X"44",X"8F",X"18",X"A0",X"2A",X"43",X"8F",
		X"7E",X"A7",X"20",X"0C",X"2A",X"41",X"8F",X"7E",X"FE",X"40",X"38",X"04",X"FE",X"C0",X"38",X"08",
		X"AF",X"21",X"40",X"8F",X"06",X"05",X"D7",X"C9",X"4F",X"3A",X"07",X"89",X"CB",X"47",X"3A",X"42",
		X"88",X"20",X"04",X"D6",X"02",X"18",X"02",X"C6",X"14",X"21",X"87",X"8A",X"47",X"3A",X"03",X"8F",
		X"3C",X"32",X"03",X"8F",X"E6",X"07",X"20",X"0D",X"78",X"C6",X"08",X"B9",X"38",X"07",X"D6",X"10",
		X"B9",X"3E",X"10",X"38",X"01",X"AF",X"77",X"78",X"B9",X"28",X"06",X"DA",X"12",X"6D",X"C3",X"0D",
		X"6D",X"CB",X"96",X"CB",X"9E",X"C9",X"3A",X"51",X"8F",X"EF",X"B8",X"6D",X"59",X"6E",X"42",X"6F",
		X"5E",X"6F",X"9D",X"6F",X"32",X"70",X"5F",X"70",X"CD",X"BC",X"0F",X"3A",X"07",X"89",X"CB",X"3F",
		X"CB",X"3F",X"FE",X"07",X"38",X"02",X"3E",X"07",X"E6",X"07",X"21",X"F3",X"70",X"CD",X"45",X"0C",
		X"ED",X"53",X"4A",X"8F",X"3E",X"40",X"32",X"48",X"8F",X"21",X"51",X"8F",X"34",X"3A",X"07",X"89",
		X"CB",X"3F",X"CB",X"3F",X"CB",X"3F",X"D0",X"21",X"C8",X"0A",X"11",X"F9",X"6D",X"06",X"60",X"1A",
		X"BE",X"C2",X"71",X"70",X"23",X"13",X"10",X"F7",X"C9",X"21",X"41",X"8D",X"35",X"20",X"03",X"CD",
		X"28",X"0A",X"CD",X"F8",X"09",X"21",X"50",X"8E",X"35",X"C0",X"36",X"02",X"2A",X"54",X"8E",X"7E",
		X"23",X"22",X"54",X"8E",X"2A",X"56",X"8E",X"77",X"11",X"E0",X"FF",X"19",X"22",X"56",X"8E",X"21",
		X"52",X"8E",X"35",X"C0",X"36",X"0D",X"21",X"50",X"8E",X"36",X"14",X"2C",X"34",X"2A",X"56",X"8E",
		X"11",X"00",X"00",X"06",X"0E",X"7E",X"83",X"5F",X"30",X"01",X"14",X"3E",X"20",X"85",X"6F",X"30",
		X"01",X"24",X"10",X"F1",X"2A",X"48",X"8F",X"7E",X"BB",X"C2",X"42",X"74",X"23",X"7E",X"BA",X"C2",
		X"EA",X"76",X"23",X"22",X"48",X"8F",X"C9",X"C6",X"01",X"CD",X"83",X"15",X"CD",X"75",X"6E",X"CD",
		X"55",X"1E",X"CD",X"D4",X"20",X"CD",X"EF",X"02",X"CD",X"DA",X"18",X"CD",X"1C",X"19",X"CD",X"04",
		X"64",X"CD",X"64",X"0E",X"C9",X"21",X"1E",X"88",X"3A",X"F0",X"8E",X"B6",X"C2",X"92",X"4C",X"CD",
		X"86",X"6E",X"CD",X"DB",X"6E",X"C9",X"21",X"48",X"8F",X"7E",X"A7",X"28",X"02",X"35",X"C9",X"3A",
		X"49",X"8F",X"CB",X"4F",X"3E",X"20",X"28",X"02",X"3E",X"2C",X"77",X"2A",X"4A",X"8F",X"7E",X"FE",
		X"FF",X"C8",X"23",X"22",X"4A",X"8F",X"47",X"DD",X"21",X"C8",X"8A",X"11",X"18",X"00",X"DD",X"19",
		X"10",X"FC",X"21",X"EA",X"8B",X"11",X"18",X"00",X"06",X"03",X"7E",X"A7",X"28",X"0B",X"19",X"10",
		X"F9",X"2A",X"4A",X"8F",X"2B",X"22",X"4A",X"8F",X"C9",X"DD",X"36",X"02",X"06",X"11",X"6A",X"39",
		X"CD",X"1E",X"38",X"CD",X"6C",X"3A",X"21",X"49",X"8F",X"34",X"C9",X"DD",X"21",X"E0",X"8A",X"11",
		X"18",X"00",X"06",X"0E",X"D9",X"CD",X"2D",X"6F",X"D9",X"DD",X"19",X"10",X"F7",X"2A",X"4A",X"8F",
		X"7E",X"FE",X"FF",X"C0",X"21",X"EA",X"8B",X"11",X"18",X"00",X"06",X"03",X"7E",X"A7",X"C0",X"19",
		X"10",X"FA",X"21",X"51",X"8F",X"34",X"23",X"11",X"35",X"06",X"FF",X"3A",X"47",X"8F",X"47",X"CB",
		X"27",X"80",X"BE",X"11",X"08",X"06",X"20",X"07",X"3E",X"04",X"32",X"51",X"8F",X"1E",X"10",X"3E",
		X"40",X"32",X"48",X"8F",X"FF",X"AF",X"21",X"90",X"8C",X"06",X"30",X"D7",X"C9",X"DD",X"7E",X"02",
		X"FE",X"02",X"CA",X"36",X"35",X"D6",X"0B",X"30",X"04",X"CD",X"06",X"40",X"C9",X"EF",X"69",X"3E",
		X"9C",X"3E",X"21",X"51",X"8F",X"34",X"23",X"7E",X"A7",X"28",X"04",X"47",X"CD",X"31",X"11",X"21",
		X"34",X"86",X"CD",X"19",X"11",X"09",X"09",X"7B",X"87",X"27",X"CD",X"19",X"11",X"C9",X"21",X"48",
		X"8F",X"7E",X"FE",X"20",X"20",X"13",X"2E",X"52",X"7E",X"A7",X"28",X"0B",X"11",X"15",X"03",X"FF",
		X"3A",X"E5",X"89",X"A7",X"C0",X"35",X"C0",X"2E",X"48",X"35",X"C0",X"36",X"60",X"3A",X"07",X"89",
		X"FE",X"03",X"C2",X"98",X"6F",X"21",X"32",X"0B",X"11",X"71",X"70",X"06",X"79",X"1A",X"BE",X"C2",
		X"F9",X"6D",X"23",X"13",X"10",X"F7",X"26",X"8F",X"2E",X"51",X"36",X"06",X"C9",X"3A",X"47",X"8F",
		X"21",X"34",X"86",X"77",X"47",X"AF",X"C6",X"05",X"10",X"FC",X"32",X"47",X"8F",X"11",X"E0",X"FF",
		X"06",X"03",X"19",X"36",X"00",X"10",X"FB",X"21",X"51",X"8F",X"34",X"2E",X"48",X"36",X"80",X"DD",
		X"21",X"C5",X"6A",X"21",X"ED",X"6F",X"06",X"44",X"DD",X"7E",X"00",X"BE",X"20",X"14",X"DD",X"2C",
		X"DD",X"7D",X"A7",X"20",X"02",X"DD",X"24",X"23",X"10",X"EE",X"CD",X"44",X"0F",X"11",X"27",X"06",
		X"FF",X"C9",X"AF",X"21",X"00",X"88",X"11",X"01",X"88",X"77",X"ED",X"B0",X"C9",X"3A",X"2D",X"89",
		X"FE",X"02",X"C0",X"3A",X"56",X"8F",X"A7",X"C0",X"3C",X"32",X"56",X"8F",X"21",X"50",X"84",X"11",
		X"00",X"00",X"7B",X"86",X"5F",X"30",X"01",X"14",X"2C",X"7D",X"E6",X"1F",X"FE",X"1B",X"20",X"03",
		X"2C",X"18",X"EF",X"FE",X"1F",X"20",X"EB",X"3E",X"12",X"85",X"6F",X"30",X"E5",X"24",X"7C",X"FE",
		X"88",X"38",X"DF",X"7B",X"FE",X"B8",X"28",X"03",X"C3",X"29",X"09",X"7A",X"FE",X"29",X"C2",X"29",
		X"38",X"C9",X"21",X"47",X"8F",X"7E",X"A7",X"C4",X"59",X"70",X"23",X"7E",X"A7",X"28",X"14",X"35",
		X"7E",X"E6",X"0F",X"A7",X"C0",X"2E",X"54",X"34",X"CB",X"46",X"11",X"A7",X"06",X"28",X"02",X"1E",
		X"27",X"FF",X"C9",X"36",X"20",X"2E",X"51",X"34",X"C9",X"35",X"11",X"15",X"03",X"FF",X"C9",X"21",
		X"48",X"8F",X"35",X"C0",X"CD",X"CF",X"0E",X"AF",X"32",X"52",X"8F",X"3E",X"06",X"32",X"0A",X"88",
		X"C9",X"21",X"BC",X"82",X"11",X"E0",X"FF",X"06",X"0A",X"7E",X"19",X"BE",X"C2",X"B3",X"08",X"10",
		X"F8",X"21",X"41",X"8D",X"35",X"20",X"03",X"CD",X"28",X"0A",X"CD",X"F8",X"09",X"21",X"50",X"8E",
		X"35",X"C0",X"36",X"01",X"2C",X"35",X"3A",X"53",X"8E",X"3D",X"21",X"AB",X"0B",X"CD",X"45",X"0C",
		X"ED",X"53",X"56",X"8E",X"21",X"53",X"8E",X"35",X"C0",X"21",X"50",X"8E",X"36",X"96",X"2C",X"AF",
		X"77",X"21",X"62",X"84",X"57",X"5F",X"0E",X"0E",X"06",X"1D",X"7B",X"86",X"30",X"01",X"14",X"5F",
		X"23",X"10",X"F7",X"7D",X"C6",X"03",X"6F",X"30",X"01",X"24",X"0D",X"20",X"EB",X"2A",X"48",X"8F",
		X"7B",X"BE",X"C2",X"B3",X"08",X"23",X"7E",X"BA",X"C2",X"E9",X"08",X"AF",X"32",X"48",X"8F",X"32",
		X"49",X"8F",X"3E",X"03",X"32",X"05",X"88",X"C3",X"00",X"0E",X"59",X"63",X"0C",X"C2",X"0B",X"62",
		X"0B",X"22",X"0B",X"03",X"71",X"13",X"71",X"26",X"71",X"3C",X"71",X"55",X"71",X"6E",X"71",X"87",
		X"71",X"A0",X"71",X"01",X"02",X"03",X"04",X"05",X"05",X"05",X"04",X"04",X"03",X"03",X"02",X"02",
		X"01",X"01",X"FF",X"01",X"01",X"02",X"02",X"03",X"03",X"04",X"04",X"05",X"05",X"06",X"06",X"06",
		X"05",X"04",X"03",X"02",X"01",X"FF",X"01",X"02",X"03",X"04",X"05",X"06",X"07",X"07",X"06",X"05",
		X"04",X"03",X"02",X"03",X"04",X"02",X"03",X"04",X"05",X"06",X"07",X"FF",X"01",X"01",X"02",X"02",
		X"03",X"03",X"04",X"04",X"05",X"05",X"06",X"06",X"07",X"07",X"08",X"08",X"08",X"07",X"06",X"05",
		X"04",X"03",X"04",X"05",X"FF",X"01",X"02",X"03",X"02",X"04",X"05",X"03",X"02",X"04",X"04",X"05",
		X"05",X"06",X"06",X"07",X"07",X"08",X"08",X"08",X"07",X"06",X"05",X"04",X"03",X"FF",X"01",X"02",
		X"03",X"04",X"05",X"06",X"07",X"08",X"08",X"07",X"06",X"05",X"04",X"03",X"02",X"01",X"01",X"02",
		X"03",X"04",X"05",X"06",X"07",X"08",X"FF",X"03",X"02",X"02",X"01",X"01",X"02",X"03",X"02",X"03",
		X"04",X"05",X"06",X"06",X"05",X"04",X"04",X"05",X"06",X"07",X"08",X"08",X"07",X"07",X"08",X"FF",
		X"01",X"02",X"03",X"04",X"05",X"06",X"07",X"08",X"08",X"08",X"07",X"07",X"06",X"06",X"05",X"05",
		X"04",X"04",X"03",X"03",X"02",X"02",X"01",X"01",X"FF",X"3A",X"38",X"8F",X"21",X"EF",X"02",X"E5",
		X"EF",X"C7",X"71",X"A0",X"72",X"21",X"74",X"CD",X"CE",X"71",X"CD",X"D4",X"20",X"C9",X"21",X"36",
		X"8F",X"7E",X"A7",X"28",X"02",X"35",X"C9",X"21",X"99",X"8A",X"3A",X"90",X"8C",X"B6",X"21",X"87",
		X"8A",X"20",X"1A",X"3A",X"5B",X"8F",X"A7",X"20",X"0F",X"3A",X"84",X"8A",X"FE",X"60",X"38",X"03",
		X"32",X"5B",X"8F",X"CB",X"96",X"CB",X"DE",X"C9",X"CB",X"D6",X"CB",X"9E",X"C9",X"3A",X"84",X"8A",
		X"FE",X"59",X"28",X"07",X"30",X"DD",X"CB",X"96",X"CB",X"DE",X"C9",X"3A",X"39",X"8F",X"A7",X"20",
		X"0A",X"3E",X"01",X"32",X"39",X"8F",X"CB",X"96",X"CB",X"9E",X"C9",X"FE",X"02",X"28",X"0B",X"3E",
		X"02",X"32",X"39",X"8F",X"3E",X"10",X"32",X"87",X"8A",X"C9",X"21",X"3E",X"8F",X"7E",X"A7",X"C2",
		X"92",X"72",X"2E",X"3B",X"34",X"7E",X"E6",X"07",X"C2",X"87",X"72",X"3A",X"96",X"8C",X"CB",X"3F",
		X"CB",X"3F",X"CB",X"3F",X"3C",X"47",X"21",X"E0",X"87",X"11",X"E0",X"FF",X"19",X"10",X"FD",X"CD",
		X"87",X"72",X"CB",X"3F",X"CB",X"3F",X"CB",X"3F",X"3C",X"47",X"23",X"10",X"FD",X"36",X"2C",X"11",
		X"00",X"FC",X"19",X"3A",X"96",X"8C",X"E6",X"06",X"FE",X"06",X"3A",X"94",X"8C",X"28",X"0C",X"E6",
		X"06",X"FE",X"02",X"28",X"03",X"36",X"00",X"C9",X"36",X"40",X"C9",X"E6",X"06",X"FE",X"02",X"28",
		X"03",X"36",X"80",X"C9",X"36",X"C0",X"C9",X"3A",X"94",X"8C",X"FE",X"D0",X"D8",X"3E",X"01",X"32",
		X"3E",X"8F",X"AF",X"32",X"87",X"8A",X"32",X"5B",X"8F",X"21",X"38",X"8F",X"34",X"23",X"77",X"C9",
		X"CD",X"D4",X"20",X"CD",X"A7",X"72",X"C9",X"21",X"3A",X"8F",X"7E",X"A7",X"20",X"04",X"CD",X"E1",
		X"72",X"C9",X"3A",X"3C",X"8F",X"A7",X"CA",X"E3",X"73",X"DD",X"21",X"E0",X"8A",X"11",X"18",X"00",
		X"3A",X"3D",X"8F",X"87",X"47",X"D9",X"CD",X"CF",X"72",X"D9",X"DD",X"19",X"10",X"F7",X"C9",X"DD",
		X"7E",X"00",X"DD",X"B6",X"01",X"0F",X"D0",X"DD",X"7E",X"02",X"EF",X"3C",X"73",X"95",X"73",X"CE",
		X"73",X"3A",X"90",X"8C",X"A7",X"C0",X"3C",X"32",X"3A",X"8F",X"21",X"3D",X"8F",X"34",X"7E",X"FE",
		X"04",X"20",X"08",X"2E",X"38",X"34",X"2E",X"36",X"36",X"20",X"C9",X"87",X"32",X"3C",X"8F",X"47",
		X"21",X"09",X"74",X"11",X"18",X"00",X"DD",X"21",X"E0",X"8A",X"DD",X"36",X"00",X"01",X"7E",X"DD",
		X"77",X"06",X"23",X"7E",X"DD",X"77",X"10",X"23",X"7E",X"DD",X"77",X"04",X"23",X"7E",X"DD",X"77",
		X"0F",X"23",X"DD",X"7D",X"CB",X"5F",X"28",X"04",X"DD",X"36",X"03",X"80",X"DD",X"36",X"05",X"80",
		X"DD",X"19",X"10",X"D6",X"78",X"21",X"38",X"8F",X"77",X"23",X"77",X"C9",X"3A",X"96",X"8C",X"CB",
		X"3F",X"CB",X"3F",X"CB",X"3F",X"DD",X"BE",X"06",X"28",X"05",X"3C",X"DD",X"BE",X"06",X"C0",X"3A",
		X"94",X"8C",X"CB",X"3F",X"CB",X"3F",X"CB",X"3F",X"C6",X"04",X"DD",X"BE",X"04",X"28",X"07",X"D8",
		X"D6",X"05",X"DD",X"BE",X"04",X"D0",X"DD",X"34",X"02",X"DD",X"7D",X"CB",X"5F",X"20",X"1B",X"11",
		X"86",X"40",X"CD",X"1E",X"38",X"DD",X"36",X"09",X"40",X"21",X"39",X"8F",X"34",X"3A",X"3D",X"8F",
		X"BE",X"C0",X"7E",X"11",X"30",X"06",X"83",X"5F",X"FF",X"C9",X"11",X"03",X"74",X"CD",X"1E",X"38",
		X"DD",X"36",X"09",X"38",X"C9",X"CD",X"06",X"40",X"DD",X"7D",X"CB",X"5F",X"20",X"18",X"DD",X"7E",
		X"03",X"DD",X"86",X"09",X"DD",X"77",X"03",X"30",X"03",X"DD",X"34",X"04",X"DD",X"7E",X"04",X"FE",
		X"1D",X"D8",X"DD",X"34",X"02",X"C9",X"DD",X"7E",X"03",X"DD",X"96",X"09",X"DD",X"77",X"03",X"30",
		X"03",X"DD",X"35",X"04",X"DD",X"7E",X"04",X"FE",X"04",X"D0",X"DD",X"34",X"02",X"C9",X"DD",X"7D",
		X"6F",X"DD",X"7C",X"67",X"AF",X"06",X"18",X"D7",X"21",X"3C",X"8F",X"35",X"C0",X"3E",X"30",X"32",
		X"36",X"8F",X"C9",X"21",X"36",X"8F",X"7E",X"A7",X"28",X"02",X"35",X"C9",X"3A",X"3D",X"8F",X"A7",
		X"28",X"06",X"11",X"B0",X"06",X"83",X"5F",X"FF",X"3E",X"18",X"32",X"36",X"8F",X"AF",X"21",X"3A",
		X"8F",X"77",X"C9",X"40",X"21",X"10",X"FF",X"03",X"74",X"0D",X"40",X"0D",X"29",X"0D",X"40",X"0B",
		X"21",X"09",X"40",X"15",X"29",X"09",X"40",X"13",X"21",X"13",X"40",X"0C",X"29",X"13",X"40",X"0A",
		X"21",X"21",X"36",X"8F",X"7E",X"A7",X"28",X"02",X"35",X"C9",X"21",X"37",X"8F",X"06",X"09",X"D7",
		X"21",X"E0",X"8A",X"06",X"48",X"D7",X"32",X"0A",X"88",X"32",X"5B",X"8F",X"3E",X"07",X"32",X"51",
		X"8E",X"C9",X"3A",X"21",X"89",X"E6",X"03",X"EF",X"4E",X"74",X"17",X"75",X"5D",X"75",X"AF",X"32",
		X"B7",X"88",X"11",X"F0",X"4A",X"21",X"E1",X"43",X"22",X"BA",X"88",X"ED",X"53",X"45",X"8F",X"21",
		X"42",X"84",X"22",X"B8",X"88",X"21",X"42",X"80",X"22",X"43",X"8F",X"21",X"21",X"89",X"34",X"21",
		X"9A",X"74",X"11",X"00",X"00",X"06",X"08",X"1A",X"BE",X"C2",X"86",X"74",X"23",X"13",X"10",X"F7",
		X"DD",X"21",X"92",X"00",X"06",X"74",X"DD",X"7E",X"00",X"BE",X"C2",X"DF",X"67",X"23",X"DD",X"2C",
		X"DD",X"7D",X"A7",X"20",X"02",X"DD",X"24",X"10",X"ED",X"C9",X"AF",X"32",X"80",X"A1",X"C3",X"92",
		X"00",X"FF",X"32",X"00",X"A0",X"31",X"00",X"90",X"32",X"00",X"88",X"06",X"08",X"C5",X"21",X"00",
		X"00",X"DD",X"21",X"79",X"00",X"11",X"00",X"00",X"4A",X"7B",X"86",X"5F",X"30",X"04",X"14",X"20",
		X"01",X"0C",X"2C",X"20",X"F4",X"24",X"7C",X"E6",X"0F",X"20",X"EE",X"32",X"00",X"A0",X"7B",X"DD",
		X"BE",X"00",X"20",X"0C",X"7A",X"DD",X"BE",X"01",X"20",X"06",X"79",X"DD",X"BE",X"02",X"28",X"02",
		X"18",X"06",X"E5",X"21",X"FF",X"8F",X"34",X"E1",X"DD",X"23",X"DD",X"23",X"DD",X"23",X"10",X"C5",
		X"3A",X"E0",X"A0",X"E6",X"0F",X"21",X"69",X"00",X"E7",X"7E",X"B7",X"18",X"16",X"57",X"E6",X"0F",
		X"5F",X"AA",X"0F",X"0F",X"0F",X"0F",X"CD",X"FA",X"00",X"7B",X"FE",X"0A",X"38",X"02",X"C6",X"07",
		X"77",X"09",X"C9",X"32",X"00",X"A0",X"CD",X"CD",X"81",X"43",X"21",X"B7",X"88",X"34",X"7E",X"FE",
		X"1C",X"C0",X"21",X"20",X"89",X"7E",X"34",X"A7",X"32",X"B7",X"88",X"C8",X"21",X"BC",X"82",X"11",
		X"00",X"00",X"0E",X"02",X"06",X"0E",X"7E",X"83",X"5F",X"30",X"01",X"14",X"7D",X"D6",X"20",X"6F",
		X"30",X"01",X"25",X"10",X"F1",X"0D",X"21",X"BC",X"86",X"20",X"E9",X"7B",X"FE",X"4F",X"C2",X"E1",
		X"43",X"15",X"C2",X"2C",X"46",X"21",X"21",X"89",X"34",X"CD",X"B2",X"0F",X"C9",X"CD",X"6D",X"75",
		X"CD",X"21",X"76",X"CD",X"13",X"6B",X"CD",X"AF",X"76",X"CD",X"EF",X"02",X"C9",X"21",X"29",X"89",
		X"7E",X"A7",X"28",X"02",X"35",X"C9",X"3A",X"2D",X"89",X"FE",X"08",X"C8",X"DD",X"21",X"E0",X"8A",
		X"FD",X"21",X"70",X"8B",X"11",X"18",X"00",X"06",X"08",X"D9",X"CD",X"95",X"75",X"D9",X"DD",X"19",
		X"FD",X"19",X"10",X"F5",X"C9",X"DD",X"7E",X"00",X"DD",X"B6",X"01",X"0F",X"D8",X"DD",X"36",X"00",
		X"01",X"AF",X"DD",X"77",X"03",X"DD",X"77",X"05",X"DD",X"36",X"04",X"15",X"DD",X"36",X"06",X"1E",
		X"3A",X"2D",X"89",X"FE",X"02",X"38",X"31",X"AF",X"FD",X"77",X"03",X"FD",X"77",X"05",X"FD",X"36",
		X"04",X"14",X"FD",X"36",X"06",X"1E",X"21",X"18",X"76",X"3A",X"22",X"89",X"E7",X"FD",X"77",X"17",
		X"21",X"57",X"56",X"CD",X"45",X"0C",X"FD",X"73",X"0C",X"FD",X"72",X"0D",X"FD",X"36",X"09",X"18",
		X"FD",X"36",X"00",X"01",X"21",X"22",X"89",X"34",X"DD",X"36",X"09",X"18",X"3A",X"2D",X"89",X"FE",
		X"02",X"38",X"02",X"3E",X"02",X"21",X"1E",X"76",X"E7",X"32",X"29",X"89",X"21",X"2D",X"89",X"34",
		X"7E",X"FE",X"03",X"11",X"DD",X"76",X"30",X"03",X"11",X"D4",X"76",X"CD",X"1E",X"38",X"3A",X"2D",
		X"89",X"87",X"87",X"FD",X"77",X"11",X"F1",X"C9",X"03",X"04",X"02",X"00",X"01",X"03",X"16",X"28",
		X"12",X"06",X"0E",X"18",X"02",X"06",X"08",X"DD",X"21",X"E0",X"8A",X"11",X"18",X"00",X"D9",X"CD",
		X"38",X"76",X"D9",X"DD",X"19",X"10",X"F7",X"C9",X"DD",X"7E",X"02",X"E6",X"03",X"EF",X"44",X"76",
		X"75",X"76",X"A6",X"76",X"DD",X"7E",X"00",X"A7",X"C8",X"CD",X"06",X"40",X"DD",X"7E",X"05",X"DD",
		X"96",X"09",X"30",X"03",X"DD",X"35",X"06",X"DD",X"77",X"05",X"DD",X"7E",X"06",X"FE",X"06",X"D0",
		X"3E",X"20",X"32",X"2E",X"89",X"11",X"18",X"00",X"06",X"0E",X"3E",X"01",X"DD",X"77",X"02",X"DD",
		X"19",X"10",X"F9",X"F1",X"C9",X"CD",X"06",X"40",X"21",X"2E",X"89",X"7E",X"A7",X"28",X"02",X"35",
		X"C9",X"3E",X"02",X"21",X"E2",X"8A",X"11",X"18",X"00",X"06",X"08",X"77",X"19",X"10",X"FC",X"AF",
		X"21",X"A2",X"8B",X"11",X"18",X"00",X"06",X"06",X"77",X"19",X"10",X"FC",X"32",X"57",X"8D",X"3E",
		X"08",X"32",X"51",X"8E",X"F1",X"C9",X"3A",X"58",X"8D",X"A7",X"C0",X"CD",X"06",X"40",X"C9",X"21",
		X"2A",X"89",X"7E",X"A7",X"28",X"02",X"35",X"C9",X"36",X"16",X"23",X"34",X"7E",X"E6",X"01",X"11",
		X"E6",X"76",X"20",X"03",X"11",X"E8",X"76",X"21",X"71",X"84",X"01",X"40",X"00",X"1A",X"77",X"13",
		X"09",X"1A",X"77",X"C9",X"45",X"0D",X"08",X"45",X"36",X"08",X"FF",X"D4",X"76",X"C0",X"03",X"08",
		X"C0",X"09",X"08",X"FF",X"DD",X"76",X"3F",X"46",X"46",X"3F",X"CD",X"F4",X"76",X"CD",X"25",X"76",
		X"CD",X"EF",X"02",X"C9",X"DD",X"21",X"A0",X"8B",X"11",X"18",X"00",X"06",X"06",X"D9",X"CD",X"07",
		X"77",X"D9",X"DD",X"19",X"10",X"F7",X"C9",X"DD",X"7E",X"00",X"DD",X"B6",X"01",X"0F",X"D0",X"DD",
		X"7E",X"02",X"E6",X"03",X"EF",X"1D",X"77",X"40",X"77",X"90",X"77",X"81",X"78",X"DD",X"35",X"11",
		X"C0",X"21",X"57",X"8D",X"7E",X"4F",X"34",X"DD",X"77",X"13",X"79",X"21",X"69",X"78",X"87",X"E7",
		X"DD",X"77",X"15",X"23",X"7E",X"DD",X"77",X"16",X"3E",X"EC",X"DD",X"77",X"0A",X"DD",X"34",X"02",
		X"CD",X"06",X"40",X"DD",X"7E",X"0A",X"ED",X"44",X"47",X"DD",X"7E",X"03",X"B8",X"30",X"03",X"DD",
		X"35",X"04",X"DD",X"86",X"0A",X"DD",X"77",X"03",X"47",X"DD",X"7E",X"04",X"E6",X"1F",X"FE",X"09",
		X"D0",X"DD",X"34",X"02",X"DD",X"36",X"11",X"18",X"CD",X"F1",X"0E",X"DD",X"7E",X"17",X"21",X"B1",
		X"41",X"CD",X"45",X"0C",X"CD",X"1E",X"38",X"11",X"B3",X"0B",X"06",X"05",X"AF",X"6F",X"67",X"1A",
		X"E6",X"1F",X"E7",X"13",X"10",X"F9",X"7D",X"84",X"C6",X"C7",X"C8",X"21",X"E9",X"89",X"34",X"C9",
		X"CD",X"06",X"40",X"DD",X"35",X"11",X"C0",X"DD",X"7E",X"13",X"21",X"21",X"78",X"CD",X"45",X"0C",
		X"DD",X"6E",X"15",X"DD",X"66",X"16",X"CD",X"0F",X"78",X"21",X"41",X"78",X"DD",X"7E",X"13",X"CD",
		X"45",X"0C",X"DD",X"6E",X"15",X"DD",X"66",X"16",X"01",X"00",X"FC",X"09",X"CD",X"0F",X"78",X"21",
		X"58",X"8D",X"7E",X"A7",X"20",X"02",X"36",X"01",X"AF",X"DD",X"77",X"00",X"DD",X"77",X"01",X"DD",
		X"77",X"02",X"DD",X"77",X"03",X"DD",X"77",X"04",X"DD",X"77",X"05",X"DD",X"77",X"06",X"DD",X"77",
		X"16",X"DD",X"7E",X"13",X"FE",X"05",X"D8",X"DD",X"36",X"01",X"01",X"DD",X"36",X"02",X"03",X"DD",
		X"36",X"11",X"80",X"21",X"BC",X"82",X"11",X"E0",X"FF",X"01",X"00",X"0A",X"7E",X"19",X"BE",X"20",
		X"74",X"81",X"4F",X"10",X"F7",X"C6",X"83",X"21",X"0E",X"78",X"BE",X"C2",X"34",X"23",X"C9",X"01",
		X"E0",X"FF",X"1A",X"77",X"13",X"23",X"1A",X"77",X"13",X"09",X"1A",X"77",X"2B",X"13",X"1A",X"77",
		X"C9",X"2D",X"78",X"31",X"78",X"31",X"78",X"35",X"78",X"39",X"78",X"3D",X"78",X"0C",X"0D",X"0C",
		X"0C",X"0C",X"0C",X"0C",X"0C",X"0E",X"0F",X"0F",X"0E",X"0C",X"3B",X"3B",X"0C",X"A4",X"A5",X"A4",
		X"A5",X"4D",X"78",X"51",X"78",X"55",X"78",X"59",X"78",X"5D",X"78",X"61",X"78",X"00",X"00",X"C0",
		X"80",X"03",X"43",X"C3",X"83",X"0D",X"4D",X"CD",X"8D",X"00",X"00",X"80",X"80",X"05",X"02",X"82",
		X"85",X"00",X"00",X"C0",X"C0",X"07",X"0D",X"0E",X"0C",X"A8",X"86",X"68",X"86",X"28",X"86",X"E8",
		X"85",X"A8",X"85",X"68",X"85",X"40",X"06",X"F0",X"FF",X"75",X"78",X"40",X"0B",X"F0",X"FF",X"75",
		X"78",X"DD",X"35",X"11",X"C0",X"FD",X"21",X"00",X"79",X"21",X"79",X"07",X"11",X"00",X"00",X"0E",
		X"09",X"06",X"20",X"7E",X"83",X"5F",X"30",X"01",X"14",X"23",X"10",X"F7",X"FD",X"7E",X"00",X"BB",
		X"C2",X"0E",X"78",X"FD",X"7E",X"01",X"BA",X"C2",X"0E",X"78",X"FD",X"7D",X"C6",X"02",X"30",X"02",
		X"FD",X"24",X"FD",X"6F",X"0D",X"20",X"DA",X"3E",X"02",X"32",X"51",X"8E",X"FD",X"21",X"48",X"85",
		X"21",X"00",X"00",X"11",X"20",X"00",X"0E",X"04",X"06",X"0C",X"FD",X"7E",X"00",X"85",X"30",X"01",
		X"24",X"6F",X"FD",X"19",X"10",X"F4",X"CB",X"41",X"20",X"08",X"11",X"E0",X"FF",X"FD",X"23",X"0D",
		X"18",X"E6",X"0D",X"28",X"07",X"11",X"FF",X"FB",X"FD",X"19",X"18",X"F6",X"7D",X"84",X"C6",X"A6",
		X"C2",X"20",X"03",X"21",X"E0",X"8A",X"AF",X"47",X"D7",X"06",X"37",X"D7",X"CD",X"C8",X"77",X"C9",
		X"B8",X"02",X"94",X"03",X"21",X"05",X"EB",X"05",X"2A",X"09",X"40",X"0A",X"41",X"0C",X"A4",X"0C",
		X"DB",X"0E",X"3A",X"06",X"88",X"A7",X"C8",X"3A",X"0D",X"88",X"A7",X"11",X"E1",X"89",X"21",X"30",
		X"8A",X"28",X"04",X"2E",X"33",X"1E",X"E2",X"1A",X"A7",X"C0",X"23",X"7E",X"2B",X"CB",X"47",X"06",
		X"3B",X"28",X"01",X"04",X"7E",X"B8",X"28",X"02",X"34",X"C9",X"36",X"00",X"23",X"34",X"7E",X"5F",
		X"E6",X"0F",X"FE",X"0A",X"C0",X"7B",X"E6",X"F0",X"C6",X"10",X"FE",X"60",X"77",X"C0",X"36",X"00",
		X"23",X"34",X"7E",X"5F",X"E6",X"0F",X"FE",X"0A",X"C0",X"7B",X"E6",X"F0",X"C6",X"10",X"77",X"C9",
		X"11",X"09",X"06",X"FF",X"DD",X"21",X"01",X"29",X"21",X"00",X"00",X"5D",X"53",X"06",X"5B",X"DD",
		X"7E",X"00",X"83",X"5F",X"30",X"01",X"14",X"4F",X"DD",X"7D",X"E6",X"01",X"20",X"06",X"79",X"85",
		X"6F",X"30",X"01",X"24",X"DD",X"23",X"10",X"E7",X"7B",X"DD",X"BE",X"00",X"C2",X"0B",X"7A",X"7A",
		X"DD",X"BE",X"01",X"C2",X"A0",X"0F",X"7D",X"DD",X"BE",X"02",X"C2",X"88",X"13",X"7C",X"DD",X"BE",
		X"03",X"C2",X"70",X"17",X"3A",X"0D",X"88",X"A7",X"DD",X"21",X"32",X"8A",X"28",X"03",X"DD",X"2E",
		X"35",X"21",X"2D",X"86",X"11",X"E0",X"FF",X"06",X"02",X"DD",X"7E",X"00",X"4F",X"E6",X"F0",X"0F",
		X"0F",X"0F",X"0F",X"77",X"19",X"79",X"E6",X"0F",X"77",X"19",X"CB",X"40",X"20",X"04",X"36",X"51",
		X"19",X"DD",X"2B",X"10",X"E4",X"DD",X"E5",X"E1",X"AF",X"06",X"03",X"D7",X"21",X"E7",X"89",X"06",
		X"07",X"7E",X"A7",X"20",X"0A",X"23",X"10",X"F9",X"C9",X"21",X"AC",X"68",X"11",X"00",X"00",X"7E",
		X"FE",X"C9",X"28",X"08",X"83",X"30",X"01",X"14",X"5F",X"23",X"18",X"F3",X"21",X"0B",X"7A",X"7B",
		X"BE",X"C2",X"D0",X"07",X"7A",X"23",X"BE",X"C2",X"85",X"1A",X"C9",X"F8",X"24",X"8D",X"7A",X"9A",
		X"7A",X"AE",X"7A",X"BB",X"7A",X"C8",X"7A",X"D5",X"7A",X"E2",X"7A",X"F2",X"7A",X"12",X"7B",X"2E",
		X"7B",X"3F",X"7B",X"53",X"7B",X"5A",X"7B",X"69",X"7B",X"7B",X"7B",X"8B",X"7B",X"C8",X"7B",X"E7",
		X"7B",X"F8",X"7B",X"08",X"7C",X"14",X"7C",X"1F",X"7C",X"2B",X"7C",X"3E",X"7C",X"4A",X"7C",X"5C",
		X"7C",X"71",X"7C",X"85",X"7C",X"8B",X"7C",X"91",X"7C",X"97",X"7C",X"A8",X"7C",X"AE",X"7C",X"B4",
		X"7C",X"BA",X"7C",X"C0",X"7C",X"C6",X"7C",X"CD",X"7C",X"DE",X"7C",X"EF",X"7C",X"FE",X"7C",X"0A",
		X"7D",X"26",X"7D",X"42",X"7D",X"53",X"7D",X"68",X"7D",X"76",X"7D",X"82",X"7D",X"98",X"7D",X"AC",
		X"7D",X"C4",X"7D",X"E2",X"7D",X"0D",X"7E",X"46",X"7E",X"56",X"7E",X"56",X"7E",X"56",X"7E",X"56",
		X"7E",X"56",X"7E",X"56",X"7E",X"56",X"7E",X"56",X"7E",X"56",X"7E",X"5A",X"7E",X"96",X"86",X"47",
		X"41",X"4D",X"45",X"40",X"40",X"4F",X"56",X"45",X"52",X"3F",X"EE",X"86",X"50",X"55",X"53",X"48",
		X"40",X"53",X"54",X"41",X"52",X"54",X"40",X"42",X"55",X"54",X"54",X"4F",X"4E",X"3F",X"94",X"86",
		X"50",X"4C",X"41",X"59",X"45",X"52",X"40",X"4F",X"4E",X"45",X"3F",X"94",X"86",X"50",X"4C",X"41",
		X"59",X"45",X"52",X"40",X"54",X"57",X"4F",X"3F",X"80",X"86",X"48",X"49",X"47",X"48",X"40",X"53",
		X"43",X"4F",X"52",X"45",X"3F",X"BF",X"87",X"40",X"43",X"52",X"45",X"44",X"49",X"54",X"40",X"40",
		X"40",X"3F",X"BF",X"87",X"40",X"46",X"52",X"45",X"45",X"40",X"50",X"4C",X"41",X"59",X"40",X"40",
		X"40",X"3F",X"38",X"87",X"4F",X"4E",X"45",X"40",X"44",X"41",X"59",X"5C",X"5C",X"5C",X"2E",X"DA",
		X"86",X"49",X"4E",X"40",X"54",X"48",X"45",X"40",X"46",X"4F",X"52",X"45",X"53",X"54",X"5C",X"5C",
		X"5C",X"3F",X"D1",X"86",X"42",X"4F",X"4E",X"55",X"53",X"40",X"50",X"4F",X"49",X"4E",X"54",X"2E",
		X"B4",X"86",X"32",X"30",X"30",X"58",X"40",X"40",X"77",X"40",X"40",X"30",X"30",X"3F",X"CA",X"86",
		X"59",X"4F",X"55",X"52",X"40",X"50",X"4C",X"41",X"59",X"40",X"54",X"49",X"4D",X"45",X"3F",X"19",
		X"87",X"4E",X"42",X"52",X"40",X"4F",X"46",X"40",X"50",X"49",X"47",X"53",X"40",X"54",X"41",X"4B",
		X"45",X"4E",X"3F",X"24",X"86",X"50",X"4C",X"41",X"59",X"3F",X"A9",X"86",X"5B",X"40",X"40",X"50",
		X"4F",X"4F",X"59",X"41",X"4E",X"40",X"40",X"5B",X"3F",X"C4",X"86",X"5B",X"40",X"40",X"43",X"48",
		X"41",X"52",X"41",X"43",X"54",X"45",X"52",X"40",X"40",X"5B",X"3F",X"A3",X"86",X"5B",X"40",X"40",
		X"50",X"4F",X"4F",X"40",X"59",X"41",X"4E",X"40",X"40",X"5B",X"3F",X"2B",X"87",X"57",X"48",X"45",
		X"4E",X"40",X"37",X"40",X"57",X"4F",X"4C",X"56",X"45",X"53",X"40",X"4A",X"4F",X"49",X"4E",X"2E",
		X"2D",X"87",X"4F",X"4E",X"40",X"54",X"48",X"45",X"40",X"43",X"4C",X"49",X"46",X"46",X"73",X"54",
		X"48",X"45",X"59",X"2E",X"2F",X"87",X"44",X"52",X"4F",X"50",X"40",X"47",X"49",X"41",X"48",X"54",
		X"40",X"52",X"4F",X"43",X"4B",X"3B",X"3B",X"3F",X"AF",X"86",X"40",X"4E",X"49",X"43",X"45",X"40",
		X"40",X"53",X"48",X"4F",X"4F",X"54",X"2E",X"D2",X"86",X"40",X"42",X"4F",X"4E",X"55",X"53",X"40",
		X"40",X"50",X"4F",X"49",X"4E",X"54",X"3F",X"BC",X"86",X"3A",X"40",X"4B",X"4F",X"4E",X"41",X"4D",
		X"49",X"40",X"40",X"31",X"39",X"38",X"32",X"3F",X"AE",X"86",X"40",X"4D",X"41",X"4D",X"41",X"73",
		X"40",X"48",X"45",X"4C",X"50",X"40",X"3B",X"3F",X"E6",X"85",X"4F",X"48",X"73",X"40",X"42",X"4F",
		X"59",X"40",X"3B",X"3F",X"56",X"87",X"40",X"4D",X"41",X"4D",X"41",X"40",X"40",X"3B",X"3F",X"19",
		X"87",X"40",X"4D",X"41",X"4D",X"41",X"40",X"40",X"3B",X"3B",X"3F",X"75",X"87",X"31",X"53",X"54",
		X"40",X"42",X"4F",X"4E",X"55",X"53",X"40",X"41",X"46",X"54",X"45",X"52",X"40",X"3F",X"75",X"85",
		X"35",X"30",X"30",X"30",X"30",X"40",X"50",X"54",X"53",X"3F",X"D1",X"86",X"4F",X"4E",X"45",X"40",
		X"50",X"4C",X"41",X"59",X"45",X"52",X"40",X"4F",X"4E",X"4C",X"59",X"3F",X"F1",X"86",X"4F",X"4E",
		X"45",X"40",X"4F",X"52",X"40",X"54",X"57",X"4F",X"40",X"50",X"4C",X"41",X"59",X"45",X"52",X"53",
		X"3F",X"04",X"87",X"5B",X"40",X"53",X"43",X"4F",X"52",X"45",X"40",X"52",X"41",X"4E",X"4B",X"49",
		X"4E",X"47",X"40",X"5B",X"3F",X"27",X"87",X"31",X"53",X"54",X"3F",X"29",X"87",X"32",X"4E",X"44",
		X"3F",X"2B",X"87",X"33",X"52",X"44",X"3F",X"2D",X"87",X"34",X"54",X"48",X"40",X"40",X"40",X"40",
		X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"3F",X"2F",X"87",X"35",X"54",X"48",X"3F",X"31",X"87",
		X"36",X"54",X"48",X"3F",X"33",X"87",X"37",X"54",X"48",X"3F",X"35",X"87",X"38",X"54",X"48",X"3F",
		X"37",X"87",X"39",X"54",X"48",X"3F",X"59",X"87",X"31",X"30",X"54",X"48",X"3F",X"BD",X"86",X"3A",
		X"40",X"4B",X"4F",X"4E",X"41",X"4D",X"49",X"40",X"40",X"31",X"39",X"38",X"32",X"3F",X"D1",X"86",
		X"40",X"42",X"4F",X"4E",X"55",X"53",X"40",X"40",X"53",X"54",X"41",X"47",X"45",X"40",X"3F",X"AC",
		X"86",X"40",X"40",X"50",X"45",X"52",X"46",X"45",X"43",X"54",X"40",X"40",X"40",X"3F",X"75",X"85",
		X"33",X"30",X"30",X"30",X"30",X"40",X"50",X"54",X"53",X"3F",X"78",X"87",X"41",X"4E",X"44",X"40",
		X"42",X"4F",X"4E",X"55",X"53",X"40",X"45",X"56",X"45",X"52",X"59",X"40",X"37",X"30",X"30",X"30",
		X"30",X"40",X"50",X"54",X"53",X"3F",X"78",X"87",X"41",X"4E",X"44",X"40",X"42",X"4F",X"4E",X"55",
		X"53",X"40",X"45",X"56",X"45",X"52",X"59",X"40",X"38",X"30",X"30",X"30",X"30",X"40",X"50",X"54",
		X"53",X"3F",X"D0",X"86",X"32",X"4E",X"44",X"40",X"50",X"48",X"41",X"53",X"45",X"40",X"47",X"45",
		X"54",X"53",X"3F",X"12",X"87",X"48",X"41",X"52",X"44",X"45",X"52",X"40",X"41",X"53",X"40",X"59",
		X"4F",X"55",X"40",X"4C",X"4F",X"53",X"45",X"3F",X"94",X"86",X"4D",X"4F",X"52",X"45",X"40",X"50",
		X"49",X"47",X"53",X"40",X"3B",X"3F",X"16",X"86",X"3F",X"44",X"49",X"46",X"46",X"49",X"43",X"55",
		X"4C",X"54",X"38",X"87",X"3F",X"49",X"4E",X"40",X"54",X"48",X"45",X"40",X"53",X"45",X"43",X"4F",
		X"4E",X"44",X"40",X"50",X"48",X"41",X"53",X"45",X"75",X"87",X"41",X"42",X"4F",X"55",X"54",X"40",
		X"31",X"30",X"40",X"53",X"45",X"43",X"4F",X"4E",X"44",X"53",X"3B",X"3F",X"92",X"86",X"40",X"4F",
		X"4E",X"45",X"40",X"57",X"4F",X"4C",X"46",X"2E",X"74",X"86",X"40",X"40",X"34",X"30",X"30",X"40",
		X"50",X"54",X"53",X"3F",X"92",X"86",X"40",X"54",X"57",X"4F",X"40",X"57",X"4F",X"4C",X"56",X"45",
		X"53",X"2E",X"74",X"86",X"40",X"40",X"34",X"30",X"30",X"83",X"38",X"30",X"30",X"40",X"50",X"54",
		X"53",X"3F",X"92",X"86",X"40",X"53",X"4F",X"4D",X"45",X"40",X"57",X"4F",X"4C",X"56",X"45",X"53",
		X"2E",X"74",X"86",X"40",X"40",X"34",X"30",X"30",X"83",X"38",X"30",X"30",X"40",X"2E",X"56",X"86",
		X"40",X"40",X"40",X"83",X"31",X"36",X"30",X"30",X"40",X"50",X"54",X"53",X"3F",X"CD",X"86",X"42",
		X"4F",X"4E",X"55",X"53",X"40",X"40",X"50",X"4F",X"49",X"4E",X"54",X"2E",X"10",X"87",X"4D",X"45",
		X"41",X"54",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"30",X"30",X"40",X"50",X"54",X"53",
		X"2E",X"12",X"87",X"57",X"4F",X"4C",X"46",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"30",
		X"30",X"40",X"50",X"54",X"53",X"3F",X"A3",X"86",X"42",X"4F",X"4E",X"55",X"53",X"40",X"40",X"53",
		X"54",X"41",X"47",X"45",X"40",X"3F",X"00",X"84",X"40",X"3F",X"89",X"86",X"44",X"4F",X"55",X"42",
		X"4C",X"45",X"2E",X"4D",X"86",X"50",X"45",X"52",X"46",X"45",X"43",X"54",X"3F",X"3A",X"88",X"89",
		X"FE",X"04",X"D8",X"3A",X"5F",X"8A",X"A7",X"C0",X"21",X"BE",X"64",X"0E",X"00",X"59",X"7E",X"2B",
		X"81",X"4F",X"30",X"01",X"1C",X"3E",X"34",X"BE",X"20",X"F4",X"7B",X"81",X"E6",X"B0",X"C8",X"21",
		X"EF",X"89",X"34",X"C9",X"21",X"D6",X"7F",X"E5",X"3A",X"2A",X"8E",X"A7",X"C0",X"3A",X"FC",X"89",
		X"A7",X"20",X"05",X"3C",X"32",X"2A",X"8E",X"C9",X"3A",X"26",X"8E",X"EF",X"B2",X"7E",X"0E",X"7F",
		X"5D",X"7F",X"21",X"65",X"85",X"22",X"27",X"8E",X"3E",X"03",X"32",X"25",X"8E",X"3A",X"FC",X"89",
		X"21",X"A0",X"03",X"22",X"2B",X"8E",X"DD",X"21",X"FD",X"8D",X"47",X"11",X"03",X"00",X"DD",X"19",
		X"10",X"FC",X"DD",X"22",X"1F",X"8E",X"3A",X"0F",X"88",X"A7",X"20",X"06",X"3A",X"0D",X"88",X"A7",
		X"20",X"05",X"21",X"11",X"88",X"18",X"03",X"21",X"12",X"88",X"22",X"21",X"8E",X"3A",X"FC",X"89",
		X"47",X"ED",X"5B",X"27",X"8E",X"13",X"13",X"10",X"FC",X"ED",X"53",X"27",X"8E",X"3E",X"11",X"12",
		X"32",X"23",X"8E",X"3E",X"01",X"32",X"26",X"8E",X"3E",X"0C",X"32",X"24",X"8E",X"C9",X"2A",X"2B",
		X"8E",X"2B",X"22",X"2B",X"8E",X"7C",X"A7",X"20",X"07",X"7D",X"A7",X"20",X"03",X"C3",X"A8",X"7F",
		X"2A",X"21",X"8E",X"CB",X"5E",X"20",X"1B",X"CB",X"56",X"28",X"32",X"21",X"24",X"8E",X"35",X"C0",
		X"3E",X"0C",X"32",X"24",X"8E",X"21",X"23",X"8E",X"34",X"7E",X"FE",X"2D",X"38",X"19",X"36",X"10",
		X"18",X"15",X"21",X"24",X"8E",X"35",X"C0",X"3E",X"0C",X"32",X"24",X"8E",X"21",X"23",X"8E",X"35",
		X"7E",X"FE",X"10",X"30",X"02",X"36",X"2C",X"ED",X"4B",X"27",X"8E",X"7E",X"02",X"2A",X"21",X"8E",
		X"7E",X"21",X"29",X"8E",X"07",X"07",X"07",X"07",X"CB",X"16",X"7E",X"E6",X"07",X"FE",X"01",X"C0",
		X"21",X"A0",X"03",X"22",X"2B",X"8E",X"3A",X"23",X"8E",X"2A",X"1F",X"8E",X"77",X"23",X"22",X"1F",
		X"8E",X"21",X"25",X"8E",X"35",X"7E",X"A7",X"32",X"25",X"8E",X"28",X"1C",X"3A",X"23",X"8E",X"2A",
		X"27",X"8E",X"77",X"01",X"E0",X"FF",X"09",X"22",X"27",X"8E",X"3E",X"11",X"77",X"3E",X"01",X"32",
		X"26",X"8E",X"3E",X"11",X"32",X"23",X"8E",X"C9",X"CD",X"CF",X"0E",X"3A",X"25",X"8E",X"A7",X"28",
		X"16",X"47",X"3E",X"10",X"2A",X"27",X"8E",X"11",X"E0",X"FF",X"DD",X"2A",X"1F",X"8E",X"77",X"DD",
		X"77",X"00",X"19",X"DD",X"23",X"10",X"F7",X"21",X"08",X"88",X"36",X"80",X"AF",X"32",X"26",X"8E",
		X"3E",X"01",X"32",X"2A",X"8E",X"C9",X"3A",X"02",X"88",X"A7",X"C8",X"21",X"0E",X"88",X"7E",X"A7",
		X"28",X"0D",X"2B",X"7E",X"A7",X"3A",X"08",X"89",X"21",X"48",X"89",X"20",X"02",X"2E",X"88",X"B6",
		X"A7",X"C0",X"3A",X"10",X"88",X"E6",X"18",X"A7",X"C8",X"CD",X"CF",X"0E",X"C3",X"78",X"0D",X"FF");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
